// Mega_JSoC.v

// Generated using ACDS version 13.1 162 at 2024.06.12.16:03:33

`timescale 1 ps / 1 ps
module Mega_JSoC (
		input  wire        clk_clk,                      //                   clk.clk
		input  wire        reset_reset_n,                //                 reset.reset_n
		output wire [12:0] sdram_controller_wire_addr,   // sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,     //                      .ba
		output wire        sdram_controller_wire_cas_n,  //                      .cas_n
		output wire        sdram_controller_wire_cke,    //                      .cke
		output wire        sdram_controller_wire_cs_n,   //                      .cs_n
		inout  wire [31:0] sdram_controller_wire_dq,     //                      .dq
		output wire [3:0]  sdram_controller_wire_dqm,    //                      .dqm
		output wire        sdram_controller_wire_ras_n,  //                      .ras_n
		output wire        sdram_controller_wire_we_n,   //                      .we_n
		input  wire        pll_areset_conduit_export,    //    pll_areset_conduit.export
		output wire        pll_locked_conduit_export,    //    pll_locked_conduit.export
		output wire        pll_phasedone_conduit_export, // pll_phasedone_conduit.export
		output wire        sdram_clk_clk                 //             sdram_clk.clk
	);

	wire         pll_c0_clk;                                                   // pll:c0 -> [cpu:clk, cpu_1b:clk, cpu_1c:clk, cpu_1d:clk, cpu_1e:clk, cpu_1f:clk, fifo_1b:wrclock, fifo_1c:wrclock, fifo_1d:wrclock, fifo_1e:wrclock, fifo_q_1:wrclock, fifo_q_2:wrclock, fifo_q_3:wrclock, fifo_q_4:wrclock, fifo_q_5:wrclock, fifo_q_6:wrclock, irq_mapper:clk, irq_mapper_001:clk, irq_mapper_002:clk, irq_mapper_003:clk, irq_mapper_004:clk, irq_mapper_005:clk, jtag_uart:clk, jtag_uart_1b:clk, jtag_uart_1c:clk, jtag_uart_1d:clk, jtag_uart_1e:clk, jtag_uart_1f:clk, mm_interconnect_0:pll_c0_clk, onchip_mem_1b:clk, onchip_mem_1c:clk, onchip_mem_1d:clk, onchip_mem_1e:clk, onchip_mem_1f:clk, rst_controller:clk, sdram_controller:clk, sys_id:clock, sysid_1b:clock, sysid_1c:clock, sysid_1d:clock, sysid_1e:clock, sysid_1f:clock, timer:clk, timer_1b:clk, timer_1c:clk, timer_1d:clk, timer_1e:clk, timer_1f:clk]
	wire         mm_interconnect_0_fifo_1d_in_waitrequest;                     // fifo_1d:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_1d_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_1d_in_writedata;                       // mm_interconnect_0:fifo_1d_in_writedata -> fifo_1d:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_1d_in_write;                           // mm_interconnect_0:fifo_1d_in_write -> fifo_1d:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo_q_6_in_waitrequest;                    // fifo_q_6:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_6_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_q_6_in_writedata;                      // mm_interconnect_0:fifo_q_6_in_writedata -> fifo_q_6:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_6_in_write;                          // mm_interconnect_0:fifo_q_6_in_write -> fifo_q_6:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo_q_4_in_waitrequest;                    // fifo_q_4:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_4_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_q_4_in_writedata;                      // mm_interconnect_0:fifo_q_4_in_writedata -> fifo_q_4:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_4_in_write;                          // mm_interconnect_0:fifo_q_4_in_write -> fifo_q_4:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_3_in_csr_writedata;                  // mm_interconnect_0:fifo_q_3_in_csr_writedata -> fifo_q_3:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_q_3_in_csr_address;                    // mm_interconnect_0:fifo_q_3_in_csr_address -> fifo_q_3:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_3_in_csr_write;                      // mm_interconnect_0:fifo_q_3_in_csr_write -> fifo_q_3:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_q_3_in_csr_read;                       // mm_interconnect_0:fifo_q_3_in_csr_read -> fifo_q_3:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_3_in_csr_readdata;                   // fifo_q_3:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_3_in_csr_readdata
	wire   [0:0] mm_interconnect_0_sys_id_control_slave_address;               // mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	wire  [31:0] mm_interconnect_0_sys_id_control_slave_readdata;              // sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	wire         cpu_1b_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_1b_instruction_master_waitrequest -> cpu_1b:i_waitrequest
	wire  [17:0] cpu_1b_instruction_master_address;                            // cpu_1b:i_address -> mm_interconnect_0:cpu_1b_instruction_master_address
	wire         cpu_1b_instruction_master_read;                               // cpu_1b:i_read -> mm_interconnect_0:cpu_1b_instruction_master_read
	wire  [31:0] cpu_1b_instruction_master_readdata;                           // mm_interconnect_0:cpu_1b_instruction_master_readdata -> cpu_1b:i_readdata
	wire         cpu_1c_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_1c_instruction_master_waitrequest -> cpu_1c:i_waitrequest
	wire  [17:0] cpu_1c_instruction_master_address;                            // cpu_1c:i_address -> mm_interconnect_0:cpu_1c_instruction_master_address
	wire         cpu_1c_instruction_master_read;                               // cpu_1c:i_read -> mm_interconnect_0:cpu_1c_instruction_master_read
	wire  [31:0] cpu_1c_instruction_master_readdata;                           // mm_interconnect_0:cpu_1c_instruction_master_readdata -> cpu_1c:i_readdata
	wire         mm_interconnect_0_cpu_1e_jtag_debug_module_waitrequest;       // cpu_1e:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_1e_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_1e_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_1e_jtag_debug_module_writedata -> cpu_1e:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_1e_jtag_debug_module_address;           // mm_interconnect_0:cpu_1e_jtag_debug_module_address -> cpu_1e:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_1e_jtag_debug_module_write;             // mm_interconnect_0:cpu_1e_jtag_debug_module_write -> cpu_1e:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_1e_jtag_debug_module_read;              // mm_interconnect_0:cpu_1e_jtag_debug_module_read -> cpu_1e:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_1e_jtag_debug_module_readdata;          // cpu_1e:jtag_debug_module_readdata -> mm_interconnect_0:cpu_1e_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_1e_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_1e_jtag_debug_module_debugaccess -> cpu_1e:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_1e_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_1e_jtag_debug_module_byteenable -> cpu_1e:jtag_debug_module_byteenable
	wire         mm_interconnect_0_fifo_q_4_out_waitrequest;                   // fifo_q_4:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_4_out_waitrequest
	wire         mm_interconnect_0_fifo_q_4_out_read;                          // mm_interconnect_0:fifo_q_4_out_read -> fifo_q_4:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_4_out_readdata;                      // fifo_q_4:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_4_out_readdata
	wire  [31:0] mm_interconnect_0_fifo_q_6_in_csr_writedata;                  // mm_interconnect_0:fifo_q_6_in_csr_writedata -> fifo_q_6:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_q_6_in_csr_address;                    // mm_interconnect_0:fifo_q_6_in_csr_address -> fifo_q_6:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_6_in_csr_write;                      // mm_interconnect_0:fifo_q_6_in_csr_write -> fifo_q_6:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_q_6_in_csr_read;                       // mm_interconnect_0:fifo_q_6_in_csr_read -> fifo_q_6:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_6_in_csr_readdata;                   // fifo_q_6:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_6_in_csr_readdata
	wire         cpu_1b_data_master_waitrequest;                               // mm_interconnect_0:cpu_1b_data_master_waitrequest -> cpu_1b:d_waitrequest
	wire  [31:0] cpu_1b_data_master_writedata;                                 // cpu_1b:d_writedata -> mm_interconnect_0:cpu_1b_data_master_writedata
	wire  [27:0] cpu_1b_data_master_address;                                   // cpu_1b:d_address -> mm_interconnect_0:cpu_1b_data_master_address
	wire         cpu_1b_data_master_write;                                     // cpu_1b:d_write -> mm_interconnect_0:cpu_1b_data_master_write
	wire         cpu_1b_data_master_read;                                      // cpu_1b:d_read -> mm_interconnect_0:cpu_1b_data_master_read
	wire  [31:0] cpu_1b_data_master_readdata;                                  // mm_interconnect_0:cpu_1b_data_master_readdata -> cpu_1b:d_readdata
	wire         cpu_1b_data_master_debugaccess;                               // cpu_1b:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_1b_data_master_debugaccess
	wire   [3:0] cpu_1b_data_master_byteenable;                                // cpu_1b:d_byteenable -> mm_interconnect_0:cpu_1b_data_master_byteenable
	wire  [31:0] mm_interconnect_0_fifo_q_5_in_csr_writedata;                  // mm_interconnect_0:fifo_q_5_in_csr_writedata -> fifo_q_5:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_q_5_in_csr_address;                    // mm_interconnect_0:fifo_q_5_in_csr_address -> fifo_q_5:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_5_in_csr_write;                      // mm_interconnect_0:fifo_q_5_in_csr_write -> fifo_q_5:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_q_5_in_csr_read;                       // mm_interconnect_0:fifo_q_5_in_csr_read -> fifo_q_5:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_5_in_csr_readdata;                   // fifo_q_5:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_5_in_csr_readdata
	wire         mm_interconnect_0_fifo_1b_out_waitrequest;                    // fifo_1b:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_1b_out_waitrequest
	wire         mm_interconnect_0_fifo_1b_out_read;                           // mm_interconnect_0:fifo_1b_out_read -> fifo_1b:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_1b_out_readdata;                       // fifo_1b:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_1b_out_readdata
	wire         cpu_1f_data_master_waitrequest;                               // mm_interconnect_0:cpu_1f_data_master_waitrequest -> cpu_1f:d_waitrequest
	wire  [31:0] cpu_1f_data_master_writedata;                                 // cpu_1f:d_writedata -> mm_interconnect_0:cpu_1f_data_master_writedata
	wire  [27:0] cpu_1f_data_master_address;                                   // cpu_1f:d_address -> mm_interconnect_0:cpu_1f_data_master_address
	wire         cpu_1f_data_master_write;                                     // cpu_1f:d_write -> mm_interconnect_0:cpu_1f_data_master_write
	wire         cpu_1f_data_master_read;                                      // cpu_1f:d_read -> mm_interconnect_0:cpu_1f_data_master_read
	wire  [31:0] cpu_1f_data_master_readdata;                                  // mm_interconnect_0:cpu_1f_data_master_readdata -> cpu_1f:d_readdata
	wire         cpu_1f_data_master_debugaccess;                               // cpu_1f:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_1f_data_master_debugaccess
	wire   [3:0] cpu_1f_data_master_byteenable;                                // cpu_1f:d_byteenable -> mm_interconnect_0:cpu_1f_data_master_byteenable
	wire         mm_interconnect_0_cpu_1d_jtag_debug_module_waitrequest;       // cpu_1d:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_1d_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_1d_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_1d_jtag_debug_module_writedata -> cpu_1d:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_1d_jtag_debug_module_address;           // mm_interconnect_0:cpu_1d_jtag_debug_module_address -> cpu_1d:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_1d_jtag_debug_module_write;             // mm_interconnect_0:cpu_1d_jtag_debug_module_write -> cpu_1d:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_1d_jtag_debug_module_read;              // mm_interconnect_0:cpu_1d_jtag_debug_module_read -> cpu_1d:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_1d_jtag_debug_module_readdata;          // cpu_1d:jtag_debug_module_readdata -> mm_interconnect_0:cpu_1d_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_1d_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_1d_jtag_debug_module_debugaccess -> cpu_1d:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_1d_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_1d_jtag_debug_module_byteenable -> cpu_1d:jtag_debug_module_byteenable
	wire         cpu_data_master_waitrequest;                                  // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                    // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [27:0] cpu_data_master_address;                                      // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                        // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                         // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                     // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                  // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                   // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         mm_interconnect_0_fifo_q_6_out_waitrequest;                   // fifo_q_6:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_6_out_waitrequest
	wire         mm_interconnect_0_fifo_q_6_out_read;                          // mm_interconnect_0:fifo_q_6_out_read -> fifo_q_6:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_6_out_readdata;                      // fifo_q_6:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_6_out_readdata
	wire  [15:0] mm_interconnect_0_timer_1b_s1_writedata;                      // mm_interconnect_0:timer_1b_s1_writedata -> timer_1b:writedata
	wire   [2:0] mm_interconnect_0_timer_1b_s1_address;                        // mm_interconnect_0:timer_1b_s1_address -> timer_1b:address
	wire         mm_interconnect_0_timer_1b_s1_chipselect;                     // mm_interconnect_0:timer_1b_s1_chipselect -> timer_1b:chipselect
	wire         mm_interconnect_0_timer_1b_s1_write;                          // mm_interconnect_0:timer_1b_s1_write -> timer_1b:write_n
	wire  [15:0] mm_interconnect_0_timer_1b_s1_readdata;                       // timer_1b:readdata -> mm_interconnect_0:timer_1b_s1_readdata
	wire  [15:0] mm_interconnect_0_timer_1c_s1_writedata;                      // mm_interconnect_0:timer_1c_s1_writedata -> timer_1c:writedata
	wire   [2:0] mm_interconnect_0_timer_1c_s1_address;                        // mm_interconnect_0:timer_1c_s1_address -> timer_1c:address
	wire         mm_interconnect_0_timer_1c_s1_chipselect;                     // mm_interconnect_0:timer_1c_s1_chipselect -> timer_1c:chipselect
	wire         mm_interconnect_0_timer_1c_s1_write;                          // mm_interconnect_0:timer_1c_s1_write -> timer_1c:write_n
	wire  [15:0] mm_interconnect_0_timer_1c_s1_readdata;                       // timer_1c:readdata -> mm_interconnect_0:timer_1c_s1_readdata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                    // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                      // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_write;                        // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire         mm_interconnect_0_pll_pll_slave_read;                         // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                     // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire         mm_interconnect_0_cpu_1c_jtag_debug_module_waitrequest;       // cpu_1c:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_1c_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_1c_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_1c_jtag_debug_module_writedata -> cpu_1c:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_1c_jtag_debug_module_address;           // mm_interconnect_0:cpu_1c_jtag_debug_module_address -> cpu_1c:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_1c_jtag_debug_module_write;             // mm_interconnect_0:cpu_1c_jtag_debug_module_write -> cpu_1c:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_1c_jtag_debug_module_read;              // mm_interconnect_0:cpu_1c_jtag_debug_module_read -> cpu_1c:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_1c_jtag_debug_module_readdata;          // cpu_1c:jtag_debug_module_readdata -> mm_interconnect_0:cpu_1c_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_1c_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_1c_jtag_debug_module_debugaccess -> cpu_1c:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_1c_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_1c_jtag_debug_module_byteenable -> cpu_1c:jtag_debug_module_byteenable
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_waitrequest; // jtag_uart_1f:av_waitrequest -> mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_writedata -> jtag_uart_1f:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_address -> jtag_uart_1f:av_address
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_chipselect -> jtag_uart_1f:av_chipselect
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_write -> jtag_uart_1f:av_write_n
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_read -> jtag_uart_1f:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_readdata;    // jtag_uart_1f:av_readdata -> mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_fifo_1c_in_csr_writedata;                   // mm_interconnect_0:fifo_1c_in_csr_writedata -> fifo_1c:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_1c_in_csr_address;                     // mm_interconnect_0:fifo_1c_in_csr_address -> fifo_1c:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_1c_in_csr_write;                       // mm_interconnect_0:fifo_1c_in_csr_write -> fifo_1c:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_1c_in_csr_read;                        // mm_interconnect_0:fifo_1c_in_csr_read -> fifo_1c:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_1c_in_csr_readdata;                    // fifo_1c:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_1c_in_csr_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;    // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;       // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_cpu_1b_jtag_debug_module_waitrequest;       // cpu_1b:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_1b_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_1b_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_1b_jtag_debug_module_writedata -> cpu_1b:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_1b_jtag_debug_module_address;           // mm_interconnect_0:cpu_1b_jtag_debug_module_address -> cpu_1b:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_1b_jtag_debug_module_write;             // mm_interconnect_0:cpu_1b_jtag_debug_module_write -> cpu_1b:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_1b_jtag_debug_module_read;              // mm_interconnect_0:cpu_1b_jtag_debug_module_read -> cpu_1b:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_1b_jtag_debug_module_readdata;          // cpu_1b:jtag_debug_module_readdata -> mm_interconnect_0:cpu_1b_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_1b_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_1b_jtag_debug_module_debugaccess -> cpu_1b:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_1b_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_1b_jtag_debug_module_byteenable -> cpu_1b:jtag_debug_module_byteenable
	wire         mm_interconnect_0_fifo_1c_in_waitrequest;                     // fifo_1c:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_1c_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_1c_in_writedata;                       // mm_interconnect_0:fifo_1c_in_writedata -> fifo_1c:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_1c_in_write;                           // mm_interconnect_0:fifo_1c_in_write -> fifo_1c:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo_1e_in_waitrequest;                     // fifo_1e:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_1e_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_1e_in_writedata;                       // mm_interconnect_0:fifo_1e_in_writedata -> fifo_1e:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_1e_in_write;                           // mm_interconnect_0:fifo_1e_in_write -> fifo_1e:avalonmm_write_slave_write
	wire   [0:0] mm_interconnect_0_sysid_1d_control_slave_address;             // mm_interconnect_0:sysid_1d_control_slave_address -> sysid_1d:address
	wire  [31:0] mm_interconnect_0_sysid_1d_control_slave_readdata;            // sysid_1d:readdata -> mm_interconnect_0:sysid_1d_control_slave_readdata
	wire         mm_interconnect_0_fifo_1d_out_waitrequest;                    // fifo_1d:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_1d_out_waitrequest
	wire         mm_interconnect_0_fifo_1d_out_read;                           // mm_interconnect_0:fifo_1d_out_read -> fifo_1d:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_1d_out_readdata;                       // fifo_1d:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_1d_out_readdata
	wire         cpu_1c_data_master_waitrequest;                               // mm_interconnect_0:cpu_1c_data_master_waitrequest -> cpu_1c:d_waitrequest
	wire  [31:0] cpu_1c_data_master_writedata;                                 // cpu_1c:d_writedata -> mm_interconnect_0:cpu_1c_data_master_writedata
	wire  [17:0] cpu_1c_data_master_address;                                   // cpu_1c:d_address -> mm_interconnect_0:cpu_1c_data_master_address
	wire         cpu_1c_data_master_write;                                     // cpu_1c:d_write -> mm_interconnect_0:cpu_1c_data_master_write
	wire         cpu_1c_data_master_read;                                      // cpu_1c:d_read -> mm_interconnect_0:cpu_1c_data_master_read
	wire  [31:0] cpu_1c_data_master_readdata;                                  // mm_interconnect_0:cpu_1c_data_master_readdata -> cpu_1c:d_readdata
	wire         cpu_1c_data_master_debugaccess;                               // cpu_1c:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_1c_data_master_debugaccess
	wire   [3:0] cpu_1c_data_master_byteenable;                                // cpu_1c:d_byteenable -> mm_interconnect_0:cpu_1c_data_master_byteenable
	wire  [31:0] mm_interconnect_0_onchip_mem_1f_s1_writedata;                 // mm_interconnect_0:onchip_mem_1f_s1_writedata -> onchip_mem_1f:writedata
	wire  [14:0] mm_interconnect_0_onchip_mem_1f_s1_address;                   // mm_interconnect_0:onchip_mem_1f_s1_address -> onchip_mem_1f:address
	wire         mm_interconnect_0_onchip_mem_1f_s1_chipselect;                // mm_interconnect_0:onchip_mem_1f_s1_chipselect -> onchip_mem_1f:chipselect
	wire         mm_interconnect_0_onchip_mem_1f_s1_clken;                     // mm_interconnect_0:onchip_mem_1f_s1_clken -> onchip_mem_1f:clken
	wire         mm_interconnect_0_onchip_mem_1f_s1_write;                     // mm_interconnect_0:onchip_mem_1f_s1_write -> onchip_mem_1f:write
	wire  [31:0] mm_interconnect_0_onchip_mem_1f_s1_readdata;                  // onchip_mem_1f:readdata -> mm_interconnect_0:onchip_mem_1f_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_mem_1f_s1_byteenable;                // mm_interconnect_0:onchip_mem_1f_s1_byteenable -> onchip_mem_1f:byteenable
	wire  [31:0] mm_interconnect_0_fifo_1e_in_csr_writedata;                   // mm_interconnect_0:fifo_1e_in_csr_writedata -> fifo_1e:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_1e_in_csr_address;                     // mm_interconnect_0:fifo_1e_in_csr_address -> fifo_1e:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_1e_in_csr_write;                       // mm_interconnect_0:fifo_1e_in_csr_write -> fifo_1e:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_1e_in_csr_read;                        // mm_interconnect_0:fifo_1e_in_csr_read -> fifo_1e:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_1e_in_csr_readdata;                    // fifo_1e:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_1e_in_csr_readdata
	wire   [0:0] mm_interconnect_0_sysid_1c_control_slave_address;             // mm_interconnect_0:sysid_1c_control_slave_address -> sysid_1c:address
	wire  [31:0] mm_interconnect_0_sysid_1c_control_slave_readdata;            // sysid_1c:readdata -> mm_interconnect_0:sysid_1c_control_slave_readdata
	wire  [31:0] mm_interconnect_0_onchip_mem_1e_s1_writedata;                 // mm_interconnect_0:onchip_mem_1e_s1_writedata -> onchip_mem_1e:writedata
	wire  [13:0] mm_interconnect_0_onchip_mem_1e_s1_address;                   // mm_interconnect_0:onchip_mem_1e_s1_address -> onchip_mem_1e:address
	wire         mm_interconnect_0_onchip_mem_1e_s1_chipselect;                // mm_interconnect_0:onchip_mem_1e_s1_chipselect -> onchip_mem_1e:chipselect
	wire         mm_interconnect_0_onchip_mem_1e_s1_clken;                     // mm_interconnect_0:onchip_mem_1e_s1_clken -> onchip_mem_1e:clken
	wire         mm_interconnect_0_onchip_mem_1e_s1_write;                     // mm_interconnect_0:onchip_mem_1e_s1_write -> onchip_mem_1e:write
	wire  [31:0] mm_interconnect_0_onchip_mem_1e_s1_readdata;                  // onchip_mem_1e:readdata -> mm_interconnect_0:onchip_mem_1e_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_mem_1e_s1_byteenable;                // mm_interconnect_0:onchip_mem_1e_s1_byteenable -> onchip_mem_1e:byteenable
	wire         cpu_1f_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_1f_instruction_master_waitrequest -> cpu_1f:i_waitrequest
	wire  [18:0] cpu_1f_instruction_master_address;                            // cpu_1f:i_address -> mm_interconnect_0:cpu_1f_instruction_master_address
	wire         cpu_1f_instruction_master_read;                               // cpu_1f:i_read -> mm_interconnect_0:cpu_1f_instruction_master_read
	wire  [31:0] cpu_1f_instruction_master_readdata;                           // mm_interconnect_0:cpu_1f_instruction_master_readdata -> cpu_1f:i_readdata
	wire  [31:0] mm_interconnect_0_onchip_mem_1d_s1_writedata;                 // mm_interconnect_0:onchip_mem_1d_s1_writedata -> onchip_mem_1d:writedata
	wire  [13:0] mm_interconnect_0_onchip_mem_1d_s1_address;                   // mm_interconnect_0:onchip_mem_1d_s1_address -> onchip_mem_1d:address
	wire         mm_interconnect_0_onchip_mem_1d_s1_chipselect;                // mm_interconnect_0:onchip_mem_1d_s1_chipselect -> onchip_mem_1d:chipselect
	wire         mm_interconnect_0_onchip_mem_1d_s1_clken;                     // mm_interconnect_0:onchip_mem_1d_s1_clken -> onchip_mem_1d:clken
	wire         mm_interconnect_0_onchip_mem_1d_s1_write;                     // mm_interconnect_0:onchip_mem_1d_s1_write -> onchip_mem_1d:write
	wire  [31:0] mm_interconnect_0_onchip_mem_1d_s1_readdata;                  // onchip_mem_1d:readdata -> mm_interconnect_0:onchip_mem_1d_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_mem_1d_s1_byteenable;                // mm_interconnect_0:onchip_mem_1d_s1_byteenable -> onchip_mem_1d:byteenable
	wire         cpu_instruction_master_waitrequest;                           // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                               // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                  // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                              // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire  [31:0] mm_interconnect_0_onchip_mem_1c_s1_writedata;                 // mm_interconnect_0:onchip_mem_1c_s1_writedata -> onchip_mem_1c:writedata
	wire  [13:0] mm_interconnect_0_onchip_mem_1c_s1_address;                   // mm_interconnect_0:onchip_mem_1c_s1_address -> onchip_mem_1c:address
	wire         mm_interconnect_0_onchip_mem_1c_s1_chipselect;                // mm_interconnect_0:onchip_mem_1c_s1_chipselect -> onchip_mem_1c:chipselect
	wire         mm_interconnect_0_onchip_mem_1c_s1_clken;                     // mm_interconnect_0:onchip_mem_1c_s1_clken -> onchip_mem_1c:clken
	wire         mm_interconnect_0_onchip_mem_1c_s1_write;                     // mm_interconnect_0:onchip_mem_1c_s1_write -> onchip_mem_1c:write
	wire  [31:0] mm_interconnect_0_onchip_mem_1c_s1_readdata;                  // onchip_mem_1c:readdata -> mm_interconnect_0:onchip_mem_1c_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_mem_1c_s1_byteenable;                // mm_interconnect_0:onchip_mem_1c_s1_byteenable -> onchip_mem_1c:byteenable
	wire   [0:0] mm_interconnect_0_sysid_1e_control_slave_address;             // mm_interconnect_0:sysid_1e_control_slave_address -> sysid_1e:address
	wire  [31:0] mm_interconnect_0_sysid_1e_control_slave_readdata;            // sysid_1e:readdata -> mm_interconnect_0:sysid_1e_control_slave_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;          // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;            // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;              // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                 // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;             // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;          // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;           // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         cpu_1e_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_1e_instruction_master_waitrequest -> cpu_1e:i_waitrequest
	wire  [17:0] cpu_1e_instruction_master_address;                            // cpu_1e:i_address -> mm_interconnect_0:cpu_1e_instruction_master_address
	wire         cpu_1e_instruction_master_read;                               // cpu_1e:i_read -> mm_interconnect_0:cpu_1e_instruction_master_read
	wire  [31:0] cpu_1e_instruction_master_readdata;                           // mm_interconnect_0:cpu_1e_instruction_master_readdata -> cpu_1e:i_readdata
	wire  [15:0] mm_interconnect_0_timer_1f_s1_writedata;                      // mm_interconnect_0:timer_1f_s1_writedata -> timer_1f:writedata
	wire   [2:0] mm_interconnect_0_timer_1f_s1_address;                        // mm_interconnect_0:timer_1f_s1_address -> timer_1f:address
	wire         mm_interconnect_0_timer_1f_s1_chipselect;                     // mm_interconnect_0:timer_1f_s1_chipselect -> timer_1f:chipselect
	wire         mm_interconnect_0_timer_1f_s1_write;                          // mm_interconnect_0:timer_1f_s1_write -> timer_1f:write_n
	wire  [15:0] mm_interconnect_0_timer_1f_s1_readdata;                       // timer_1f:readdata -> mm_interconnect_0:timer_1f_s1_readdata
	wire   [0:0] mm_interconnect_0_sysid_1b_control_slave_address;             // mm_interconnect_0:sysid_1b_control_slave_address -> sysid_1b:address
	wire  [31:0] mm_interconnect_0_sysid_1b_control_slave_readdata;            // sysid_1b:readdata -> mm_interconnect_0:sysid_1b_control_slave_readdata
	wire  [31:0] mm_interconnect_0_fifo_q_1_in_csr_writedata;                  // mm_interconnect_0:fifo_q_1_in_csr_writedata -> fifo_q_1:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_q_1_in_csr_address;                    // mm_interconnect_0:fifo_q_1_in_csr_address -> fifo_q_1:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_1_in_csr_write;                      // mm_interconnect_0:fifo_q_1_in_csr_write -> fifo_q_1:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_q_1_in_csr_read;                       // mm_interconnect_0:fifo_q_1_in_csr_read -> fifo_q_1:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_1_in_csr_readdata;                   // fifo_q_1:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_1_in_csr_readdata
	wire  [31:0] mm_interconnect_0_fifo_1b_in_csr_writedata;                   // mm_interconnect_0:fifo_1b_in_csr_writedata -> fifo_1b:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_1b_in_csr_address;                     // mm_interconnect_0:fifo_1b_in_csr_address -> fifo_1b:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_1b_in_csr_write;                       // mm_interconnect_0:fifo_1b_in_csr_write -> fifo_1b:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_1b_in_csr_read;                        // mm_interconnect_0:fifo_1b_in_csr_read -> fifo_1b:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_1b_in_csr_readdata;                    // fifo_1b:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_1b_in_csr_readdata
	wire         mm_interconnect_0_fifo_q_2_out_waitrequest;                   // fifo_q_2:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_2_out_waitrequest
	wire         mm_interconnect_0_fifo_q_2_out_read;                          // mm_interconnect_0:fifo_q_2_out_read -> fifo_q_2:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_2_out_readdata;                      // fifo_q_2:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_2_out_readdata
	wire         mm_interconnect_0_fifo_q_5_in_waitrequest;                    // fifo_q_5:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_5_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_q_5_in_writedata;                      // mm_interconnect_0:fifo_q_5_in_writedata -> fifo_q_5:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_5_in_write;                          // mm_interconnect_0:fifo_q_5_in_write -> fifo_q_5:avalonmm_write_slave_write
	wire         mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_waitrequest; // jtag_uart_1d:av_waitrequest -> mm_interconnect_0:jtag_uart_1d_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1d_avalon_jtag_slave_writedata -> jtag_uart_1d:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1d_avalon_jtag_slave_address -> jtag_uart_1d:av_address
	wire         mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1d_avalon_jtag_slave_chipselect -> jtag_uart_1d:av_chipselect
	wire         mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1d_avalon_jtag_slave_write -> jtag_uart_1d:av_write_n
	wire         mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1d_avalon_jtag_slave_read -> jtag_uart_1d:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_readdata;    // jtag_uart_1d:av_readdata -> mm_interconnect_0:jtag_uart_1d_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_waitrequest; // jtag_uart_1e:av_waitrequest -> mm_interconnect_0:jtag_uart_1e_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1e_avalon_jtag_slave_writedata -> jtag_uart_1e:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1e_avalon_jtag_slave_address -> jtag_uart_1e:av_address
	wire         mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1e_avalon_jtag_slave_chipselect -> jtag_uart_1e:av_chipselect
	wire         mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1e_avalon_jtag_slave_write -> jtag_uart_1e:av_write_n
	wire         mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1e_avalon_jtag_slave_read -> jtag_uart_1e:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_readdata;    // jtag_uart_1e:av_readdata -> mm_interconnect_0:jtag_uart_1e_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_onchip_mem_1b_s1_writedata;                 // mm_interconnect_0:onchip_mem_1b_s1_writedata -> onchip_mem_1b:writedata
	wire  [13:0] mm_interconnect_0_onchip_mem_1b_s1_address;                   // mm_interconnect_0:onchip_mem_1b_s1_address -> onchip_mem_1b:address
	wire         mm_interconnect_0_onchip_mem_1b_s1_chipselect;                // mm_interconnect_0:onchip_mem_1b_s1_chipselect -> onchip_mem_1b:chipselect
	wire         mm_interconnect_0_onchip_mem_1b_s1_clken;                     // mm_interconnect_0:onchip_mem_1b_s1_clken -> onchip_mem_1b:clken
	wire         mm_interconnect_0_onchip_mem_1b_s1_write;                     // mm_interconnect_0:onchip_mem_1b_s1_write -> onchip_mem_1b:write
	wire  [31:0] mm_interconnect_0_onchip_mem_1b_s1_readdata;                  // onchip_mem_1b:readdata -> mm_interconnect_0:onchip_mem_1b_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_mem_1b_s1_byteenable;                // mm_interconnect_0:onchip_mem_1b_s1_byteenable -> onchip_mem_1b:byteenable
	wire         mm_interconnect_0_fifo_q_1_out_waitrequest;                   // fifo_q_1:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_1_out_waitrequest
	wire         mm_interconnect_0_fifo_q_1_out_read;                          // mm_interconnect_0:fifo_q_1_out_read -> fifo_q_1:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_1_out_readdata;                      // fifo_q_1:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_1_out_readdata
	wire         mm_interconnect_0_cpu_1f_jtag_debug_module_waitrequest;       // cpu_1f:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_1f_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_1f_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_1f_jtag_debug_module_writedata -> cpu_1f:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_1f_jtag_debug_module_address;           // mm_interconnect_0:cpu_1f_jtag_debug_module_address -> cpu_1f:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_1f_jtag_debug_module_write;             // mm_interconnect_0:cpu_1f_jtag_debug_module_write -> cpu_1f:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_1f_jtag_debug_module_read;              // mm_interconnect_0:cpu_1f_jtag_debug_module_read -> cpu_1f:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_1f_jtag_debug_module_readdata;          // cpu_1f:jtag_debug_module_readdata -> mm_interconnect_0:cpu_1f_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_1f_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_1f_jtag_debug_module_debugaccess -> cpu_1f:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_1f_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_1f_jtag_debug_module_byteenable -> cpu_1f:jtag_debug_module_byteenable
	wire         mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_waitrequest; // jtag_uart_1c:av_waitrequest -> mm_interconnect_0:jtag_uart_1c_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1c_avalon_jtag_slave_writedata -> jtag_uart_1c:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1c_avalon_jtag_slave_address -> jtag_uart_1c:av_address
	wire         mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1c_avalon_jtag_slave_chipselect -> jtag_uart_1c:av_chipselect
	wire         mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1c_avalon_jtag_slave_write -> jtag_uart_1c:av_write_n
	wire         mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1c_avalon_jtag_slave_read -> jtag_uart_1c:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_readdata;    // jtag_uart_1c:av_readdata -> mm_interconnect_0:jtag_uart_1c_avalon_jtag_slave_readdata
	wire         cpu_1e_data_master_waitrequest;                               // mm_interconnect_0:cpu_1e_data_master_waitrequest -> cpu_1e:d_waitrequest
	wire  [31:0] cpu_1e_data_master_writedata;                                 // cpu_1e:d_writedata -> mm_interconnect_0:cpu_1e_data_master_writedata
	wire  [27:0] cpu_1e_data_master_address;                                   // cpu_1e:d_address -> mm_interconnect_0:cpu_1e_data_master_address
	wire         cpu_1e_data_master_write;                                     // cpu_1e:d_write -> mm_interconnect_0:cpu_1e_data_master_write
	wire         cpu_1e_data_master_read;                                      // cpu_1e:d_read -> mm_interconnect_0:cpu_1e_data_master_read
	wire  [31:0] cpu_1e_data_master_readdata;                                  // mm_interconnect_0:cpu_1e_data_master_readdata -> cpu_1e:d_readdata
	wire         cpu_1e_data_master_debugaccess;                               // cpu_1e:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_1e_data_master_debugaccess
	wire   [3:0] cpu_1e_data_master_byteenable;                                // cpu_1e:d_byteenable -> mm_interconnect_0:cpu_1e_data_master_byteenable
	wire   [0:0] mm_interconnect_0_sysid_1f_control_slave_address;             // mm_interconnect_0:sysid_1f_control_slave_address -> sysid_1f:address
	wire  [31:0] mm_interconnect_0_sysid_1f_control_slave_readdata;            // sysid_1f:readdata -> mm_interconnect_0:sysid_1f_control_slave_readdata
	wire         mm_interconnect_0_fifo_1b_in_waitrequest;                     // fifo_1b:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_1b_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_1b_in_writedata;                       // mm_interconnect_0:fifo_1b_in_writedata -> fifo_1b:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_1b_in_write;                           // mm_interconnect_0:fifo_1b_in_write -> fifo_1b:avalonmm_write_slave_write
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;            // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;              // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;                // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;             // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire         mm_interconnect_0_sdram_controller_s1_write;                  // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire         mm_interconnect_0_sdram_controller_s1_read;                   // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;               // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;          // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;             // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         cpu_1d_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_1d_instruction_master_waitrequest -> cpu_1d:i_waitrequest
	wire  [17:0] cpu_1d_instruction_master_address;                            // cpu_1d:i_address -> mm_interconnect_0:cpu_1d_instruction_master_address
	wire         cpu_1d_instruction_master_read;                               // cpu_1d:i_read -> mm_interconnect_0:cpu_1d_instruction_master_read
	wire  [31:0] cpu_1d_instruction_master_readdata;                           // mm_interconnect_0:cpu_1d_instruction_master_readdata -> cpu_1d:i_readdata
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                         // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                           // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_chipselect;                        // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_0_timer_s1_write;                             // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                          // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire  [31:0] mm_interconnect_0_fifo_q_2_in_csr_writedata;                  // mm_interconnect_0:fifo_q_2_in_csr_writedata -> fifo_q_2:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_q_2_in_csr_address;                    // mm_interconnect_0:fifo_q_2_in_csr_address -> fifo_q_2:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_2_in_csr_write;                      // mm_interconnect_0:fifo_q_2_in_csr_write -> fifo_q_2:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_q_2_in_csr_read;                       // mm_interconnect_0:fifo_q_2_in_csr_read -> fifo_q_2:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_2_in_csr_readdata;                   // fifo_q_2:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_2_in_csr_readdata
	wire         mm_interconnect_0_fifo_q_1_in_waitrequest;                    // fifo_q_1:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_1_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_q_1_in_writedata;                      // mm_interconnect_0:fifo_q_1_in_writedata -> fifo_q_1:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_1_in_write;                          // mm_interconnect_0:fifo_q_1_in_write -> fifo_q_1:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_4_in_csr_writedata;                  // mm_interconnect_0:fifo_q_4_in_csr_writedata -> fifo_q_4:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_q_4_in_csr_address;                    // mm_interconnect_0:fifo_q_4_in_csr_address -> fifo_q_4:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_4_in_csr_write;                      // mm_interconnect_0:fifo_q_4_in_csr_write -> fifo_q_4:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_q_4_in_csr_read;                       // mm_interconnect_0:fifo_q_4_in_csr_read -> fifo_q_4:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_4_in_csr_readdata;                   // fifo_q_4:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_4_in_csr_readdata
	wire         mm_interconnect_0_fifo_q_2_in_waitrequest;                    // fifo_q_2:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_2_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_q_2_in_writedata;                      // mm_interconnect_0:fifo_q_2_in_writedata -> fifo_q_2:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_2_in_write;                          // mm_interconnect_0:fifo_q_2_in_write -> fifo_q_2:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo_1e_out_waitrequest;                    // fifo_1e:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_1e_out_waitrequest
	wire         mm_interconnect_0_fifo_1e_out_read;                           // mm_interconnect_0:fifo_1e_out_read -> fifo_1e:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_1e_out_readdata;                       // fifo_1e:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_1e_out_readdata
	wire         mm_interconnect_0_fifo_q_3_in_waitrequest;                    // fifo_q_3:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_3_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_q_3_in_writedata;                      // mm_interconnect_0:fifo_q_3_in_writedata -> fifo_q_3:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_3_in_write;                          // mm_interconnect_0:fifo_q_3_in_write -> fifo_q_3:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_1d_in_csr_writedata;                   // mm_interconnect_0:fifo_1d_in_csr_writedata -> fifo_1d:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_1d_in_csr_address;                     // mm_interconnect_0:fifo_1d_in_csr_address -> fifo_1d:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_1d_in_csr_write;                       // mm_interconnect_0:fifo_1d_in_csr_write -> fifo_1d:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_1d_in_csr_read;                        // mm_interconnect_0:fifo_1d_in_csr_read -> fifo_1d:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_1d_in_csr_readdata;                    // fifo_1d:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_1d_in_csr_readdata
	wire  [15:0] mm_interconnect_0_timer_1d_s1_writedata;                      // mm_interconnect_0:timer_1d_s1_writedata -> timer_1d:writedata
	wire   [2:0] mm_interconnect_0_timer_1d_s1_address;                        // mm_interconnect_0:timer_1d_s1_address -> timer_1d:address
	wire         mm_interconnect_0_timer_1d_s1_chipselect;                     // mm_interconnect_0:timer_1d_s1_chipselect -> timer_1d:chipselect
	wire         mm_interconnect_0_timer_1d_s1_write;                          // mm_interconnect_0:timer_1d_s1_write -> timer_1d:write_n
	wire  [15:0] mm_interconnect_0_timer_1d_s1_readdata;                       // timer_1d:readdata -> mm_interconnect_0:timer_1d_s1_readdata
	wire  [15:0] mm_interconnect_0_timer_1e_s1_writedata;                      // mm_interconnect_0:timer_1e_s1_writedata -> timer_1e:writedata
	wire   [2:0] mm_interconnect_0_timer_1e_s1_address;                        // mm_interconnect_0:timer_1e_s1_address -> timer_1e:address
	wire         mm_interconnect_0_timer_1e_s1_chipselect;                     // mm_interconnect_0:timer_1e_s1_chipselect -> timer_1e:chipselect
	wire         mm_interconnect_0_timer_1e_s1_write;                          // mm_interconnect_0:timer_1e_s1_write -> timer_1e:write_n
	wire  [15:0] mm_interconnect_0_timer_1e_s1_readdata;                       // timer_1e:readdata -> mm_interconnect_0:timer_1e_s1_readdata
	wire         mm_interconnect_0_fifo_q_3_out_waitrequest;                   // fifo_q_3:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_3_out_waitrequest
	wire         mm_interconnect_0_fifo_q_3_out_read;                          // mm_interconnect_0:fifo_q_3_out_read -> fifo_q_3:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_3_out_readdata;                      // fifo_q_3:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_3_out_readdata
	wire         cpu_1d_data_master_waitrequest;                               // mm_interconnect_0:cpu_1d_data_master_waitrequest -> cpu_1d:d_waitrequest
	wire  [31:0] cpu_1d_data_master_writedata;                                 // cpu_1d:d_writedata -> mm_interconnect_0:cpu_1d_data_master_writedata
	wire  [27:0] cpu_1d_data_master_address;                                   // cpu_1d:d_address -> mm_interconnect_0:cpu_1d_data_master_address
	wire         cpu_1d_data_master_write;                                     // cpu_1d:d_write -> mm_interconnect_0:cpu_1d_data_master_write
	wire         cpu_1d_data_master_read;                                      // cpu_1d:d_read -> mm_interconnect_0:cpu_1d_data_master_read
	wire  [31:0] cpu_1d_data_master_readdata;                                  // mm_interconnect_0:cpu_1d_data_master_readdata -> cpu_1d:d_readdata
	wire         cpu_1d_data_master_debugaccess;                               // cpu_1d:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_1d_data_master_debugaccess
	wire   [3:0] cpu_1d_data_master_byteenable;                                // cpu_1d:d_byteenable -> mm_interconnect_0:cpu_1d_data_master_byteenable
	wire         mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_waitrequest; // jtag_uart_1b:av_waitrequest -> mm_interconnect_0:jtag_uart_1b_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1b_avalon_jtag_slave_writedata -> jtag_uart_1b:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1b_avalon_jtag_slave_address -> jtag_uart_1b:av_address
	wire         mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1b_avalon_jtag_slave_chipselect -> jtag_uart_1b:av_chipselect
	wire         mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1b_avalon_jtag_slave_write -> jtag_uart_1b:av_write_n
	wire         mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1b_avalon_jtag_slave_read -> jtag_uart_1b:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_readdata;    // jtag_uart_1b:av_readdata -> mm_interconnect_0:jtag_uart_1b_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_fifo_1c_out_waitrequest;                    // fifo_1c:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_1c_out_waitrequest
	wire         mm_interconnect_0_fifo_1c_out_read;                           // mm_interconnect_0:fifo_1c_out_read -> fifo_1c:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_1c_out_readdata;                       // fifo_1c:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_1c_out_readdata
	wire         mm_interconnect_0_fifo_q_5_out_waitrequest;                   // fifo_q_5:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_5_out_waitrequest
	wire         mm_interconnect_0_fifo_q_5_out_read;                          // mm_interconnect_0:fifo_q_5_out_read -> fifo_q_5:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_5_out_readdata;                      // fifo_q_5:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_5_out_readdata
	wire         irq_mapper_receiver0_irq;                                     // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_d_irq_irq;                                                // irq_mapper:sender_irq -> cpu:d_irq
	wire         irq_mapper_001_receiver0_irq;                                 // timer_1b:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                 // jtag_uart_1b:av_irq -> irq_mapper_001:receiver1_irq
	wire  [31:0] cpu_1b_d_irq_irq;                                             // irq_mapper_001:sender_irq -> cpu_1b:d_irq
	wire         irq_mapper_002_receiver0_irq;                                 // timer_1c:irq -> irq_mapper_002:receiver0_irq
	wire         irq_mapper_002_receiver1_irq;                                 // jtag_uart_1c:av_irq -> irq_mapper_002:receiver1_irq
	wire  [31:0] cpu_1c_d_irq_irq;                                             // irq_mapper_002:sender_irq -> cpu_1c:d_irq
	wire         irq_mapper_003_receiver0_irq;                                 // timer_1d:irq -> irq_mapper_003:receiver0_irq
	wire         irq_mapper_003_receiver1_irq;                                 // jtag_uart_1d:av_irq -> irq_mapper_003:receiver1_irq
	wire  [31:0] cpu_1d_d_irq_irq;                                             // irq_mapper_003:sender_irq -> cpu_1d:d_irq
	wire         irq_mapper_004_receiver0_irq;                                 // timer_1e:irq -> irq_mapper_004:receiver0_irq
	wire         irq_mapper_004_receiver1_irq;                                 // jtag_uart_1e:av_irq -> irq_mapper_004:receiver1_irq
	wire  [31:0] cpu_1e_d_irq_irq;                                             // irq_mapper_004:sender_irq -> cpu_1e:d_irq
	wire         irq_mapper_005_receiver0_irq;                                 // timer_1f:irq -> irq_mapper_005:receiver0_irq
	wire         irq_mapper_005_receiver1_irq;                                 // jtag_uart_1f:av_irq -> irq_mapper_005:receiver1_irq
	wire  [31:0] cpu_1f_d_irq_irq;                                             // irq_mapper_005:sender_irq -> cpu_1f:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [cpu:reset_n, cpu_1b:reset_n, cpu_1c:reset_n, cpu_1d:reset_n, cpu_1e:reset_n, cpu_1f:reset_n, fifo_1b:reset_n, fifo_1c:reset_n, fifo_1d:reset_n, fifo_1e:reset_n, fifo_q_1:reset_n, fifo_q_2:reset_n, fifo_q_3:reset_n, fifo_q_4:reset_n, fifo_q_5:reset_n, fifo_q_6:reset_n, irq_mapper:reset, irq_mapper_001:reset, irq_mapper_002:reset, irq_mapper_003:reset, irq_mapper_004:reset, irq_mapper_005:reset, jtag_uart:rst_n, jtag_uart_1b:rst_n, jtag_uart_1c:rst_n, jtag_uart_1d:rst_n, jtag_uart_1e:rst_n, jtag_uart_1f:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_mem_1b:reset, onchip_mem_1c:reset, onchip_mem_1d:reset, onchip_mem_1e:reset, onchip_mem_1f:reset, rst_translator:in_reset, sdram_controller:reset_n, sys_id:reset_n, sysid_1b:reset_n, sysid_1c:reset_n, sysid_1d:reset_n, sysid_1e:reset_n, sysid_1f:reset_n, timer:reset_n, timer_1b:reset_n, timer_1c:reset_n, timer_1d:reset_n, timer_1e:reset_n, timer_1f:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [cpu:reset_req, cpu_1b:reset_req, cpu_1c:reset_req, cpu_1d:reset_req, cpu_1e:reset_req, cpu_1f:reset_req, onchip_mem_1b:reset_req, onchip_mem_1c:reset_req, onchip_mem_1d:reset_req, onchip_mem_1e:reset_req, onchip_mem_1f:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                            // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         cpu_1b_jtag_debug_module_reset_reset;                         // cpu_1b:jtag_debug_module_resetrequest -> [rst_controller:reset_in2, rst_controller_001:reset_in2]
	wire         cpu_1c_jtag_debug_module_reset_reset;                         // cpu_1c:jtag_debug_module_resetrequest -> [rst_controller:reset_in3, rst_controller_001:reset_in3]
	wire         cpu_1d_jtag_debug_module_reset_reset;                         // cpu_1d:jtag_debug_module_resetrequest -> [rst_controller:reset_in4, rst_controller_001:reset_in4]
	wire         cpu_1e_jtag_debug_module_reset_reset;                         // cpu_1e:jtag_debug_module_resetrequest -> [rst_controller:reset_in5, rst_controller_001:reset_in5]
	wire         cpu_1f_jtag_debug_module_reset_reset;                         // cpu_1f:jtag_debug_module_resetrequest -> [rst_controller:reset_in6, rst_controller_001:reset_in6]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	Mega_JSoC_timer timer (
		.clk        (pll_c0_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	Mega_JSoC_sys_id sys_id (
		.clock    (pll_c0_clk),                                      //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //              .address
	);

	Mega_JSoC_jtag_uart jtag_uart (
		.clk            (pll_c0_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	Mega_JSoC_cpu cpu (
		.clk                                   (pll_c0_clk),                                          //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	Mega_JSoC_sdram_controller sdram_controller (
		.clk            (pll_c0_clk),                                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                           //      .export
	);

	Mega_JSoC_pll pll (
		.clk       (clk_clk),                                   //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),        // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                             //                    c1.clk
		.areset    (pll_areset_conduit_export),                 //        areset_conduit.export
		.locked    (pll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (pll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	Mega_JSoC_cpu_1b cpu_1b (
		.clk                                   (pll_c0_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                        //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                             (cpu_1b_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_1b_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_1b_data_master_read),                                //                          .read
		.d_readdata                            (cpu_1b_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_1b_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_1b_data_master_write),                               //                          .write
		.d_writedata                           (cpu_1b_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_1b_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_1b_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_1b_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_1b_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_1b_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_1b_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_1b_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_1b_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_1b_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_1b_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_1b_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_1b_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_1b_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_1b_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_1b_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                        // custom_instruction_master.readra
	);

	Mega_JSoC_timer timer_1b (
		.clk        (pll_c0_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_1b_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1b_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1b_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1b_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1b_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver0_irq)              //   irq.irq
	);

	Mega_JSoC_onchip_mem_1b onchip_mem_1b (
		.clk        (pll_c0_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_mem_1b_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_mem_1b_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_mem_1b_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_mem_1b_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_mem_1b_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_mem_1b_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_mem_1b_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	Mega_JSoC_jtag_uart jtag_uart_1b (
		.clk            (pll_c0_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver1_irq)                                  //               irq.irq
	);

	Mega_JSoC_sysid_1b sysid_1b (
		.clock    (pll_c0_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_1b_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_1b_control_slave_address)   //              .address
	);

	Mega_JSoC_fifo_1b fifo_1b (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),            // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_1b_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_1b_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_1b_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_1b_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_1b_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_1b_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_1b_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_1b_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_1b_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_1b_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_1b_in_csr_readdata)   //         .readdata
	);

	Mega_JSoC_cpu_1c cpu_1c (
		.clk                                   (pll_c0_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                        //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                             (cpu_1c_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_1c_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_1c_data_master_read),                                //                          .read
		.d_readdata                            (cpu_1c_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_1c_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_1c_data_master_write),                               //                          .write
		.d_writedata                           (cpu_1c_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_1c_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_1c_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_1c_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_1c_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_1c_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_1c_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_1c_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_1c_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_1c_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_1c_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_1c_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_1c_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_1c_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_1c_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_1c_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                        // custom_instruction_master.readra
	);

	Mega_JSoC_timer timer_1c (
		.clk        (pll_c0_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_1c_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1c_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1c_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1c_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1c_s1_write),     //      .write_n
		.irq        (irq_mapper_002_receiver0_irq)              //   irq.irq
	);

	Mega_JSoC_onchip_mem_1c onchip_mem_1c (
		.clk        (pll_c0_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_mem_1c_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_mem_1c_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_mem_1c_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_mem_1c_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_mem_1c_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_mem_1c_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_mem_1c_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	Mega_JSoC_jtag_uart jtag_uart_1c (
		.clk            (pll_c0_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_002_receiver1_irq)                                  //               irq.irq
	);

	Mega_JSoC_sysid_1c sysid_1c (
		.clock    (pll_c0_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_1c_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_1c_control_slave_address)   //              .address
	);

	Mega_JSoC_fifo_1b fifo_1c (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),            // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_1c_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_1c_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_1c_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_1c_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_1c_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_1c_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_1c_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_1c_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_1c_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_1c_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_1c_in_csr_readdata)   //         .readdata
	);

	Mega_JSoC_cpu_1d cpu_1d (
		.clk                                   (pll_c0_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                        //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                             (cpu_1d_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_1d_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_1d_data_master_read),                                //                          .read
		.d_readdata                            (cpu_1d_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_1d_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_1d_data_master_write),                               //                          .write
		.d_writedata                           (cpu_1d_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_1d_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_1d_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_1d_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_1d_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_1d_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_1d_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_1d_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_1d_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_1d_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_1d_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_1d_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_1d_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_1d_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_1d_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_1d_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                        // custom_instruction_master.readra
	);

	Mega_JSoC_timer timer_1d (
		.clk        (pll_c0_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_1d_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1d_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1d_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1d_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1d_s1_write),     //      .write_n
		.irq        (irq_mapper_003_receiver0_irq)              //   irq.irq
	);

	Mega_JSoC_onchip_mem_1d onchip_mem_1d (
		.clk        (pll_c0_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_mem_1d_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_mem_1d_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_mem_1d_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_mem_1d_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_mem_1d_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_mem_1d_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_mem_1d_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	Mega_JSoC_jtag_uart jtag_uart_1d (
		.clk            (pll_c0_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_003_receiver1_irq)                                  //               irq.irq
	);

	Mega_JSoC_sysid_1d sysid_1d (
		.clock    (pll_c0_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_1d_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_1d_control_slave_address)   //              .address
	);

	Mega_JSoC_fifo_1b fifo_1d (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),            // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_1d_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_1d_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_1d_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_1d_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_1d_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_1d_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_1d_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_1d_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_1d_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_1d_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_1d_in_csr_readdata)   //         .readdata
	);

	Mega_JSoC_cpu_1e cpu_1e (
		.clk                                   (pll_c0_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                        //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                             (cpu_1e_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_1e_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_1e_data_master_read),                                //                          .read
		.d_readdata                            (cpu_1e_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_1e_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_1e_data_master_write),                               //                          .write
		.d_writedata                           (cpu_1e_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_1e_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_1e_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_1e_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_1e_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_1e_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_1e_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_1e_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_1e_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_1e_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_1e_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_1e_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_1e_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_1e_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_1e_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_1e_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                        // custom_instruction_master.readra
	);

	Mega_JSoC_timer timer_1e (
		.clk        (pll_c0_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_1e_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1e_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1e_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1e_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1e_s1_write),     //      .write_n
		.irq        (irq_mapper_004_receiver0_irq)              //   irq.irq
	);

	Mega_JSoC_onchip_mem_1e onchip_mem_1e (
		.clk        (pll_c0_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_mem_1e_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_mem_1e_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_mem_1e_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_mem_1e_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_mem_1e_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_mem_1e_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_mem_1e_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	Mega_JSoC_jtag_uart jtag_uart_1e (
		.clk            (pll_c0_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_004_receiver1_irq)                                  //               irq.irq
	);

	Mega_JSoC_sysid_1e sysid_1e (
		.clock    (pll_c0_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_1e_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_1e_control_slave_address)   //              .address
	);

	Mega_JSoC_fifo_1b fifo_1e (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),            // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_1e_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_1e_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_1e_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_1e_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_1e_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_1e_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_1e_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_1e_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_1e_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_1e_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_1e_in_csr_readdata)   //         .readdata
	);

	Mega_JSoC_cpu_1f cpu_1f (
		.clk                                   (pll_c0_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                        //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                             (cpu_1f_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_1f_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_1f_data_master_read),                                //                          .read
		.d_readdata                            (cpu_1f_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_1f_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_1f_data_master_write),                               //                          .write
		.d_writedata                           (cpu_1f_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_1f_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_1f_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_1f_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_1f_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_1f_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_1f_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_1f_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_1f_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_1f_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_1f_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_1f_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_1f_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_1f_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_1f_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_1f_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                        // custom_instruction_master.readra
	);

	Mega_JSoC_timer timer_1f (
		.clk        (pll_c0_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_1f_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1f_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1f_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1f_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1f_s1_write),     //      .write_n
		.irq        (irq_mapper_005_receiver0_irq)              //   irq.irq
	);

	Mega_JSoC_onchip_mem_1f onchip_mem_1f (
		.clk        (pll_c0_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_mem_1f_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_mem_1f_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_mem_1f_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_mem_1f_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_mem_1f_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_mem_1f_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_mem_1f_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	Mega_JSoC_jtag_uart jtag_uart_1f (
		.clk            (pll_c0_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_005_receiver1_irq)                                  //               irq.irq
	);

	Mega_JSoC_sysid_1f sysid_1f (
		.clock    (pll_c0_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_1f_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_1f_control_slave_address)   //              .address
	);

	Mega_JSoC_fifo_q_1 fifo_q_1 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),             // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_1_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_1_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_1_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_1_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_1_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_1_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_1_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_1_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_1_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_1_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_1_in_csr_readdata)   //         .readdata
	);

	Mega_JSoC_fifo_q_1 fifo_q_2 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),             // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_2_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_2_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_2_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_2_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_2_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_2_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_2_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_2_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_2_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_2_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_2_in_csr_readdata)   //         .readdata
	);

	Mega_JSoC_fifo_q_1 fifo_q_3 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),             // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_3_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_3_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_3_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_3_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_3_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_3_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_3_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_3_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_3_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_3_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_3_in_csr_readdata)   //         .readdata
	);

	Mega_JSoC_fifo_1b fifo_q_4 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),             // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_4_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_4_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_4_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_4_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_4_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_4_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_4_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_4_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_4_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_4_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_4_in_csr_readdata)   //         .readdata
	);

	Mega_JSoC_fifo_1b fifo_q_5 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),             // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_5_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_5_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_5_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_5_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_5_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_5_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_5_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_5_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_5_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_5_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_5_in_csr_readdata)   //         .readdata
	);

	Mega_JSoC_fifo_1b fifo_q_6 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),             // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_6_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_6_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_6_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_6_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_6_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_6_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_6_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_6_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_6_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_6_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_6_in_csr_readdata)   //         .readdata
	);

	Mega_JSoC_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                         (clk_clk),                                                      //                                       clock_clk.clk
		.pll_c0_clk                                            (pll_c0_clk),                                                   //                                          pll_c0.clk
		.cpu_reset_n_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                               //               cpu_reset_n_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                           // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                               (cpu_data_master_address),                                      //                                 cpu_data_master.address
		.cpu_data_master_waitrequest                           (cpu_data_master_waitrequest),                                  //                                                .waitrequest
		.cpu_data_master_byteenable                            (cpu_data_master_byteenable),                                   //                                                .byteenable
		.cpu_data_master_read                                  (cpu_data_master_read),                                         //                                                .read
		.cpu_data_master_readdata                              (cpu_data_master_readdata),                                     //                                                .readdata
		.cpu_data_master_write                                 (cpu_data_master_write),                                        //                                                .write
		.cpu_data_master_writedata                             (cpu_data_master_writedata),                                    //                                                .writedata
		.cpu_data_master_debugaccess                           (cpu_data_master_debugaccess),                                  //                                                .debugaccess
		.cpu_instruction_master_address                        (cpu_instruction_master_address),                               //                          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                    (cpu_instruction_master_waitrequest),                           //                                                .waitrequest
		.cpu_instruction_master_read                           (cpu_instruction_master_read),                                  //                                                .read
		.cpu_instruction_master_readdata                       (cpu_instruction_master_readdata),                              //                                                .readdata
		.cpu_1b_data_master_address                            (cpu_1b_data_master_address),                                   //                              cpu_1b_data_master.address
		.cpu_1b_data_master_waitrequest                        (cpu_1b_data_master_waitrequest),                               //                                                .waitrequest
		.cpu_1b_data_master_byteenable                         (cpu_1b_data_master_byteenable),                                //                                                .byteenable
		.cpu_1b_data_master_read                               (cpu_1b_data_master_read),                                      //                                                .read
		.cpu_1b_data_master_readdata                           (cpu_1b_data_master_readdata),                                  //                                                .readdata
		.cpu_1b_data_master_write                              (cpu_1b_data_master_write),                                     //                                                .write
		.cpu_1b_data_master_writedata                          (cpu_1b_data_master_writedata),                                 //                                                .writedata
		.cpu_1b_data_master_debugaccess                        (cpu_1b_data_master_debugaccess),                               //                                                .debugaccess
		.cpu_1b_instruction_master_address                     (cpu_1b_instruction_master_address),                            //                       cpu_1b_instruction_master.address
		.cpu_1b_instruction_master_waitrequest                 (cpu_1b_instruction_master_waitrequest),                        //                                                .waitrequest
		.cpu_1b_instruction_master_read                        (cpu_1b_instruction_master_read),                               //                                                .read
		.cpu_1b_instruction_master_readdata                    (cpu_1b_instruction_master_readdata),                           //                                                .readdata
		.cpu_1c_data_master_address                            (cpu_1c_data_master_address),                                   //                              cpu_1c_data_master.address
		.cpu_1c_data_master_waitrequest                        (cpu_1c_data_master_waitrequest),                               //                                                .waitrequest
		.cpu_1c_data_master_byteenable                         (cpu_1c_data_master_byteenable),                                //                                                .byteenable
		.cpu_1c_data_master_read                               (cpu_1c_data_master_read),                                      //                                                .read
		.cpu_1c_data_master_readdata                           (cpu_1c_data_master_readdata),                                  //                                                .readdata
		.cpu_1c_data_master_write                              (cpu_1c_data_master_write),                                     //                                                .write
		.cpu_1c_data_master_writedata                          (cpu_1c_data_master_writedata),                                 //                                                .writedata
		.cpu_1c_data_master_debugaccess                        (cpu_1c_data_master_debugaccess),                               //                                                .debugaccess
		.cpu_1c_instruction_master_address                     (cpu_1c_instruction_master_address),                            //                       cpu_1c_instruction_master.address
		.cpu_1c_instruction_master_waitrequest                 (cpu_1c_instruction_master_waitrequest),                        //                                                .waitrequest
		.cpu_1c_instruction_master_read                        (cpu_1c_instruction_master_read),                               //                                                .read
		.cpu_1c_instruction_master_readdata                    (cpu_1c_instruction_master_readdata),                           //                                                .readdata
		.cpu_1d_data_master_address                            (cpu_1d_data_master_address),                                   //                              cpu_1d_data_master.address
		.cpu_1d_data_master_waitrequest                        (cpu_1d_data_master_waitrequest),                               //                                                .waitrequest
		.cpu_1d_data_master_byteenable                         (cpu_1d_data_master_byteenable),                                //                                                .byteenable
		.cpu_1d_data_master_read                               (cpu_1d_data_master_read),                                      //                                                .read
		.cpu_1d_data_master_readdata                           (cpu_1d_data_master_readdata),                                  //                                                .readdata
		.cpu_1d_data_master_write                              (cpu_1d_data_master_write),                                     //                                                .write
		.cpu_1d_data_master_writedata                          (cpu_1d_data_master_writedata),                                 //                                                .writedata
		.cpu_1d_data_master_debugaccess                        (cpu_1d_data_master_debugaccess),                               //                                                .debugaccess
		.cpu_1d_instruction_master_address                     (cpu_1d_instruction_master_address),                            //                       cpu_1d_instruction_master.address
		.cpu_1d_instruction_master_waitrequest                 (cpu_1d_instruction_master_waitrequest),                        //                                                .waitrequest
		.cpu_1d_instruction_master_read                        (cpu_1d_instruction_master_read),                               //                                                .read
		.cpu_1d_instruction_master_readdata                    (cpu_1d_instruction_master_readdata),                           //                                                .readdata
		.cpu_1e_data_master_address                            (cpu_1e_data_master_address),                                   //                              cpu_1e_data_master.address
		.cpu_1e_data_master_waitrequest                        (cpu_1e_data_master_waitrequest),                               //                                                .waitrequest
		.cpu_1e_data_master_byteenable                         (cpu_1e_data_master_byteenable),                                //                                                .byteenable
		.cpu_1e_data_master_read                               (cpu_1e_data_master_read),                                      //                                                .read
		.cpu_1e_data_master_readdata                           (cpu_1e_data_master_readdata),                                  //                                                .readdata
		.cpu_1e_data_master_write                              (cpu_1e_data_master_write),                                     //                                                .write
		.cpu_1e_data_master_writedata                          (cpu_1e_data_master_writedata),                                 //                                                .writedata
		.cpu_1e_data_master_debugaccess                        (cpu_1e_data_master_debugaccess),                               //                                                .debugaccess
		.cpu_1e_instruction_master_address                     (cpu_1e_instruction_master_address),                            //                       cpu_1e_instruction_master.address
		.cpu_1e_instruction_master_waitrequest                 (cpu_1e_instruction_master_waitrequest),                        //                                                .waitrequest
		.cpu_1e_instruction_master_read                        (cpu_1e_instruction_master_read),                               //                                                .read
		.cpu_1e_instruction_master_readdata                    (cpu_1e_instruction_master_readdata),                           //                                                .readdata
		.cpu_1f_data_master_address                            (cpu_1f_data_master_address),                                   //                              cpu_1f_data_master.address
		.cpu_1f_data_master_waitrequest                        (cpu_1f_data_master_waitrequest),                               //                                                .waitrequest
		.cpu_1f_data_master_byteenable                         (cpu_1f_data_master_byteenable),                                //                                                .byteenable
		.cpu_1f_data_master_read                               (cpu_1f_data_master_read),                                      //                                                .read
		.cpu_1f_data_master_readdata                           (cpu_1f_data_master_readdata),                                  //                                                .readdata
		.cpu_1f_data_master_write                              (cpu_1f_data_master_write),                                     //                                                .write
		.cpu_1f_data_master_writedata                          (cpu_1f_data_master_writedata),                                 //                                                .writedata
		.cpu_1f_data_master_debugaccess                        (cpu_1f_data_master_debugaccess),                               //                                                .debugaccess
		.cpu_1f_instruction_master_address                     (cpu_1f_instruction_master_address),                            //                       cpu_1f_instruction_master.address
		.cpu_1f_instruction_master_waitrequest                 (cpu_1f_instruction_master_waitrequest),                        //                                                .waitrequest
		.cpu_1f_instruction_master_read                        (cpu_1f_instruction_master_read),                               //                                                .read
		.cpu_1f_instruction_master_readdata                    (cpu_1f_instruction_master_readdata),                           //                                                .readdata
		.cpu_jtag_debug_module_address                         (mm_interconnect_0_cpu_jtag_debug_module_address),              //                           cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                           (mm_interconnect_0_cpu_jtag_debug_module_write),                //                                                .write
		.cpu_jtag_debug_module_read                            (mm_interconnect_0_cpu_jtag_debug_module_read),                 //                                                .read
		.cpu_jtag_debug_module_readdata                        (mm_interconnect_0_cpu_jtag_debug_module_readdata),             //                                                .readdata
		.cpu_jtag_debug_module_writedata                       (mm_interconnect_0_cpu_jtag_debug_module_writedata),            //                                                .writedata
		.cpu_jtag_debug_module_byteenable                      (mm_interconnect_0_cpu_jtag_debug_module_byteenable),           //                                                .byteenable
		.cpu_jtag_debug_module_waitrequest                     (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),          //                                                .waitrequest
		.cpu_jtag_debug_module_debugaccess                     (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),          //                                                .debugaccess
		.cpu_1b_jtag_debug_module_address                      (mm_interconnect_0_cpu_1b_jtag_debug_module_address),           //                        cpu_1b_jtag_debug_module.address
		.cpu_1b_jtag_debug_module_write                        (mm_interconnect_0_cpu_1b_jtag_debug_module_write),             //                                                .write
		.cpu_1b_jtag_debug_module_read                         (mm_interconnect_0_cpu_1b_jtag_debug_module_read),              //                                                .read
		.cpu_1b_jtag_debug_module_readdata                     (mm_interconnect_0_cpu_1b_jtag_debug_module_readdata),          //                                                .readdata
		.cpu_1b_jtag_debug_module_writedata                    (mm_interconnect_0_cpu_1b_jtag_debug_module_writedata),         //                                                .writedata
		.cpu_1b_jtag_debug_module_byteenable                   (mm_interconnect_0_cpu_1b_jtag_debug_module_byteenable),        //                                                .byteenable
		.cpu_1b_jtag_debug_module_waitrequest                  (mm_interconnect_0_cpu_1b_jtag_debug_module_waitrequest),       //                                                .waitrequest
		.cpu_1b_jtag_debug_module_debugaccess                  (mm_interconnect_0_cpu_1b_jtag_debug_module_debugaccess),       //                                                .debugaccess
		.cpu_1c_jtag_debug_module_address                      (mm_interconnect_0_cpu_1c_jtag_debug_module_address),           //                        cpu_1c_jtag_debug_module.address
		.cpu_1c_jtag_debug_module_write                        (mm_interconnect_0_cpu_1c_jtag_debug_module_write),             //                                                .write
		.cpu_1c_jtag_debug_module_read                         (mm_interconnect_0_cpu_1c_jtag_debug_module_read),              //                                                .read
		.cpu_1c_jtag_debug_module_readdata                     (mm_interconnect_0_cpu_1c_jtag_debug_module_readdata),          //                                                .readdata
		.cpu_1c_jtag_debug_module_writedata                    (mm_interconnect_0_cpu_1c_jtag_debug_module_writedata),         //                                                .writedata
		.cpu_1c_jtag_debug_module_byteenable                   (mm_interconnect_0_cpu_1c_jtag_debug_module_byteenable),        //                                                .byteenable
		.cpu_1c_jtag_debug_module_waitrequest                  (mm_interconnect_0_cpu_1c_jtag_debug_module_waitrequest),       //                                                .waitrequest
		.cpu_1c_jtag_debug_module_debugaccess                  (mm_interconnect_0_cpu_1c_jtag_debug_module_debugaccess),       //                                                .debugaccess
		.cpu_1d_jtag_debug_module_address                      (mm_interconnect_0_cpu_1d_jtag_debug_module_address),           //                        cpu_1d_jtag_debug_module.address
		.cpu_1d_jtag_debug_module_write                        (mm_interconnect_0_cpu_1d_jtag_debug_module_write),             //                                                .write
		.cpu_1d_jtag_debug_module_read                         (mm_interconnect_0_cpu_1d_jtag_debug_module_read),              //                                                .read
		.cpu_1d_jtag_debug_module_readdata                     (mm_interconnect_0_cpu_1d_jtag_debug_module_readdata),          //                                                .readdata
		.cpu_1d_jtag_debug_module_writedata                    (mm_interconnect_0_cpu_1d_jtag_debug_module_writedata),         //                                                .writedata
		.cpu_1d_jtag_debug_module_byteenable                   (mm_interconnect_0_cpu_1d_jtag_debug_module_byteenable),        //                                                .byteenable
		.cpu_1d_jtag_debug_module_waitrequest                  (mm_interconnect_0_cpu_1d_jtag_debug_module_waitrequest),       //                                                .waitrequest
		.cpu_1d_jtag_debug_module_debugaccess                  (mm_interconnect_0_cpu_1d_jtag_debug_module_debugaccess),       //                                                .debugaccess
		.cpu_1e_jtag_debug_module_address                      (mm_interconnect_0_cpu_1e_jtag_debug_module_address),           //                        cpu_1e_jtag_debug_module.address
		.cpu_1e_jtag_debug_module_write                        (mm_interconnect_0_cpu_1e_jtag_debug_module_write),             //                                                .write
		.cpu_1e_jtag_debug_module_read                         (mm_interconnect_0_cpu_1e_jtag_debug_module_read),              //                                                .read
		.cpu_1e_jtag_debug_module_readdata                     (mm_interconnect_0_cpu_1e_jtag_debug_module_readdata),          //                                                .readdata
		.cpu_1e_jtag_debug_module_writedata                    (mm_interconnect_0_cpu_1e_jtag_debug_module_writedata),         //                                                .writedata
		.cpu_1e_jtag_debug_module_byteenable                   (mm_interconnect_0_cpu_1e_jtag_debug_module_byteenable),        //                                                .byteenable
		.cpu_1e_jtag_debug_module_waitrequest                  (mm_interconnect_0_cpu_1e_jtag_debug_module_waitrequest),       //                                                .waitrequest
		.cpu_1e_jtag_debug_module_debugaccess                  (mm_interconnect_0_cpu_1e_jtag_debug_module_debugaccess),       //                                                .debugaccess
		.cpu_1f_jtag_debug_module_address                      (mm_interconnect_0_cpu_1f_jtag_debug_module_address),           //                        cpu_1f_jtag_debug_module.address
		.cpu_1f_jtag_debug_module_write                        (mm_interconnect_0_cpu_1f_jtag_debug_module_write),             //                                                .write
		.cpu_1f_jtag_debug_module_read                         (mm_interconnect_0_cpu_1f_jtag_debug_module_read),              //                                                .read
		.cpu_1f_jtag_debug_module_readdata                     (mm_interconnect_0_cpu_1f_jtag_debug_module_readdata),          //                                                .readdata
		.cpu_1f_jtag_debug_module_writedata                    (mm_interconnect_0_cpu_1f_jtag_debug_module_writedata),         //                                                .writedata
		.cpu_1f_jtag_debug_module_byteenable                   (mm_interconnect_0_cpu_1f_jtag_debug_module_byteenable),        //                                                .byteenable
		.cpu_1f_jtag_debug_module_waitrequest                  (mm_interconnect_0_cpu_1f_jtag_debug_module_waitrequest),       //                                                .waitrequest
		.cpu_1f_jtag_debug_module_debugaccess                  (mm_interconnect_0_cpu_1f_jtag_debug_module_debugaccess),       //                                                .debugaccess
		.fifo_1b_in_write                                      (mm_interconnect_0_fifo_1b_in_write),                           //                                      fifo_1b_in.write
		.fifo_1b_in_writedata                                  (mm_interconnect_0_fifo_1b_in_writedata),                       //                                                .writedata
		.fifo_1b_in_waitrequest                                (mm_interconnect_0_fifo_1b_in_waitrequest),                     //                                                .waitrequest
		.fifo_1b_in_csr_address                                (mm_interconnect_0_fifo_1b_in_csr_address),                     //                                  fifo_1b_in_csr.address
		.fifo_1b_in_csr_write                                  (mm_interconnect_0_fifo_1b_in_csr_write),                       //                                                .write
		.fifo_1b_in_csr_read                                   (mm_interconnect_0_fifo_1b_in_csr_read),                        //                                                .read
		.fifo_1b_in_csr_readdata                               (mm_interconnect_0_fifo_1b_in_csr_readdata),                    //                                                .readdata
		.fifo_1b_in_csr_writedata                              (mm_interconnect_0_fifo_1b_in_csr_writedata),                   //                                                .writedata
		.fifo_1b_out_read                                      (mm_interconnect_0_fifo_1b_out_read),                           //                                     fifo_1b_out.read
		.fifo_1b_out_readdata                                  (mm_interconnect_0_fifo_1b_out_readdata),                       //                                                .readdata
		.fifo_1b_out_waitrequest                               (mm_interconnect_0_fifo_1b_out_waitrequest),                    //                                                .waitrequest
		.fifo_1c_in_write                                      (mm_interconnect_0_fifo_1c_in_write),                           //                                      fifo_1c_in.write
		.fifo_1c_in_writedata                                  (mm_interconnect_0_fifo_1c_in_writedata),                       //                                                .writedata
		.fifo_1c_in_waitrequest                                (mm_interconnect_0_fifo_1c_in_waitrequest),                     //                                                .waitrequest
		.fifo_1c_in_csr_address                                (mm_interconnect_0_fifo_1c_in_csr_address),                     //                                  fifo_1c_in_csr.address
		.fifo_1c_in_csr_write                                  (mm_interconnect_0_fifo_1c_in_csr_write),                       //                                                .write
		.fifo_1c_in_csr_read                                   (mm_interconnect_0_fifo_1c_in_csr_read),                        //                                                .read
		.fifo_1c_in_csr_readdata                               (mm_interconnect_0_fifo_1c_in_csr_readdata),                    //                                                .readdata
		.fifo_1c_in_csr_writedata                              (mm_interconnect_0_fifo_1c_in_csr_writedata),                   //                                                .writedata
		.fifo_1c_out_read                                      (mm_interconnect_0_fifo_1c_out_read),                           //                                     fifo_1c_out.read
		.fifo_1c_out_readdata                                  (mm_interconnect_0_fifo_1c_out_readdata),                       //                                                .readdata
		.fifo_1c_out_waitrequest                               (mm_interconnect_0_fifo_1c_out_waitrequest),                    //                                                .waitrequest
		.fifo_1d_in_write                                      (mm_interconnect_0_fifo_1d_in_write),                           //                                      fifo_1d_in.write
		.fifo_1d_in_writedata                                  (mm_interconnect_0_fifo_1d_in_writedata),                       //                                                .writedata
		.fifo_1d_in_waitrequest                                (mm_interconnect_0_fifo_1d_in_waitrequest),                     //                                                .waitrequest
		.fifo_1d_in_csr_address                                (mm_interconnect_0_fifo_1d_in_csr_address),                     //                                  fifo_1d_in_csr.address
		.fifo_1d_in_csr_write                                  (mm_interconnect_0_fifo_1d_in_csr_write),                       //                                                .write
		.fifo_1d_in_csr_read                                   (mm_interconnect_0_fifo_1d_in_csr_read),                        //                                                .read
		.fifo_1d_in_csr_readdata                               (mm_interconnect_0_fifo_1d_in_csr_readdata),                    //                                                .readdata
		.fifo_1d_in_csr_writedata                              (mm_interconnect_0_fifo_1d_in_csr_writedata),                   //                                                .writedata
		.fifo_1d_out_read                                      (mm_interconnect_0_fifo_1d_out_read),                           //                                     fifo_1d_out.read
		.fifo_1d_out_readdata                                  (mm_interconnect_0_fifo_1d_out_readdata),                       //                                                .readdata
		.fifo_1d_out_waitrequest                               (mm_interconnect_0_fifo_1d_out_waitrequest),                    //                                                .waitrequest
		.fifo_1e_in_write                                      (mm_interconnect_0_fifo_1e_in_write),                           //                                      fifo_1e_in.write
		.fifo_1e_in_writedata                                  (mm_interconnect_0_fifo_1e_in_writedata),                       //                                                .writedata
		.fifo_1e_in_waitrequest                                (mm_interconnect_0_fifo_1e_in_waitrequest),                     //                                                .waitrequest
		.fifo_1e_in_csr_address                                (mm_interconnect_0_fifo_1e_in_csr_address),                     //                                  fifo_1e_in_csr.address
		.fifo_1e_in_csr_write                                  (mm_interconnect_0_fifo_1e_in_csr_write),                       //                                                .write
		.fifo_1e_in_csr_read                                   (mm_interconnect_0_fifo_1e_in_csr_read),                        //                                                .read
		.fifo_1e_in_csr_readdata                               (mm_interconnect_0_fifo_1e_in_csr_readdata),                    //                                                .readdata
		.fifo_1e_in_csr_writedata                              (mm_interconnect_0_fifo_1e_in_csr_writedata),                   //                                                .writedata
		.fifo_1e_out_read                                      (mm_interconnect_0_fifo_1e_out_read),                           //                                     fifo_1e_out.read
		.fifo_1e_out_readdata                                  (mm_interconnect_0_fifo_1e_out_readdata),                       //                                                .readdata
		.fifo_1e_out_waitrequest                               (mm_interconnect_0_fifo_1e_out_waitrequest),                    //                                                .waitrequest
		.fifo_q_1_in_write                                     (mm_interconnect_0_fifo_q_1_in_write),                          //                                     fifo_q_1_in.write
		.fifo_q_1_in_writedata                                 (mm_interconnect_0_fifo_q_1_in_writedata),                      //                                                .writedata
		.fifo_q_1_in_waitrequest                               (mm_interconnect_0_fifo_q_1_in_waitrequest),                    //                                                .waitrequest
		.fifo_q_1_in_csr_address                               (mm_interconnect_0_fifo_q_1_in_csr_address),                    //                                 fifo_q_1_in_csr.address
		.fifo_q_1_in_csr_write                                 (mm_interconnect_0_fifo_q_1_in_csr_write),                      //                                                .write
		.fifo_q_1_in_csr_read                                  (mm_interconnect_0_fifo_q_1_in_csr_read),                       //                                                .read
		.fifo_q_1_in_csr_readdata                              (mm_interconnect_0_fifo_q_1_in_csr_readdata),                   //                                                .readdata
		.fifo_q_1_in_csr_writedata                             (mm_interconnect_0_fifo_q_1_in_csr_writedata),                  //                                                .writedata
		.fifo_q_1_out_read                                     (mm_interconnect_0_fifo_q_1_out_read),                          //                                    fifo_q_1_out.read
		.fifo_q_1_out_readdata                                 (mm_interconnect_0_fifo_q_1_out_readdata),                      //                                                .readdata
		.fifo_q_1_out_waitrequest                              (mm_interconnect_0_fifo_q_1_out_waitrequest),                   //                                                .waitrequest
		.fifo_q_2_in_write                                     (mm_interconnect_0_fifo_q_2_in_write),                          //                                     fifo_q_2_in.write
		.fifo_q_2_in_writedata                                 (mm_interconnect_0_fifo_q_2_in_writedata),                      //                                                .writedata
		.fifo_q_2_in_waitrequest                               (mm_interconnect_0_fifo_q_2_in_waitrequest),                    //                                                .waitrequest
		.fifo_q_2_in_csr_address                               (mm_interconnect_0_fifo_q_2_in_csr_address),                    //                                 fifo_q_2_in_csr.address
		.fifo_q_2_in_csr_write                                 (mm_interconnect_0_fifo_q_2_in_csr_write),                      //                                                .write
		.fifo_q_2_in_csr_read                                  (mm_interconnect_0_fifo_q_2_in_csr_read),                       //                                                .read
		.fifo_q_2_in_csr_readdata                              (mm_interconnect_0_fifo_q_2_in_csr_readdata),                   //                                                .readdata
		.fifo_q_2_in_csr_writedata                             (mm_interconnect_0_fifo_q_2_in_csr_writedata),                  //                                                .writedata
		.fifo_q_2_out_read                                     (mm_interconnect_0_fifo_q_2_out_read),                          //                                    fifo_q_2_out.read
		.fifo_q_2_out_readdata                                 (mm_interconnect_0_fifo_q_2_out_readdata),                      //                                                .readdata
		.fifo_q_2_out_waitrequest                              (mm_interconnect_0_fifo_q_2_out_waitrequest),                   //                                                .waitrequest
		.fifo_q_3_in_write                                     (mm_interconnect_0_fifo_q_3_in_write),                          //                                     fifo_q_3_in.write
		.fifo_q_3_in_writedata                                 (mm_interconnect_0_fifo_q_3_in_writedata),                      //                                                .writedata
		.fifo_q_3_in_waitrequest                               (mm_interconnect_0_fifo_q_3_in_waitrequest),                    //                                                .waitrequest
		.fifo_q_3_in_csr_address                               (mm_interconnect_0_fifo_q_3_in_csr_address),                    //                                 fifo_q_3_in_csr.address
		.fifo_q_3_in_csr_write                                 (mm_interconnect_0_fifo_q_3_in_csr_write),                      //                                                .write
		.fifo_q_3_in_csr_read                                  (mm_interconnect_0_fifo_q_3_in_csr_read),                       //                                                .read
		.fifo_q_3_in_csr_readdata                              (mm_interconnect_0_fifo_q_3_in_csr_readdata),                   //                                                .readdata
		.fifo_q_3_in_csr_writedata                             (mm_interconnect_0_fifo_q_3_in_csr_writedata),                  //                                                .writedata
		.fifo_q_3_out_read                                     (mm_interconnect_0_fifo_q_3_out_read),                          //                                    fifo_q_3_out.read
		.fifo_q_3_out_readdata                                 (mm_interconnect_0_fifo_q_3_out_readdata),                      //                                                .readdata
		.fifo_q_3_out_waitrequest                              (mm_interconnect_0_fifo_q_3_out_waitrequest),                   //                                                .waitrequest
		.fifo_q_4_in_write                                     (mm_interconnect_0_fifo_q_4_in_write),                          //                                     fifo_q_4_in.write
		.fifo_q_4_in_writedata                                 (mm_interconnect_0_fifo_q_4_in_writedata),                      //                                                .writedata
		.fifo_q_4_in_waitrequest                               (mm_interconnect_0_fifo_q_4_in_waitrequest),                    //                                                .waitrequest
		.fifo_q_4_in_csr_address                               (mm_interconnect_0_fifo_q_4_in_csr_address),                    //                                 fifo_q_4_in_csr.address
		.fifo_q_4_in_csr_write                                 (mm_interconnect_0_fifo_q_4_in_csr_write),                      //                                                .write
		.fifo_q_4_in_csr_read                                  (mm_interconnect_0_fifo_q_4_in_csr_read),                       //                                                .read
		.fifo_q_4_in_csr_readdata                              (mm_interconnect_0_fifo_q_4_in_csr_readdata),                   //                                                .readdata
		.fifo_q_4_in_csr_writedata                             (mm_interconnect_0_fifo_q_4_in_csr_writedata),                  //                                                .writedata
		.fifo_q_4_out_read                                     (mm_interconnect_0_fifo_q_4_out_read),                          //                                    fifo_q_4_out.read
		.fifo_q_4_out_readdata                                 (mm_interconnect_0_fifo_q_4_out_readdata),                      //                                                .readdata
		.fifo_q_4_out_waitrequest                              (mm_interconnect_0_fifo_q_4_out_waitrequest),                   //                                                .waitrequest
		.fifo_q_5_in_write                                     (mm_interconnect_0_fifo_q_5_in_write),                          //                                     fifo_q_5_in.write
		.fifo_q_5_in_writedata                                 (mm_interconnect_0_fifo_q_5_in_writedata),                      //                                                .writedata
		.fifo_q_5_in_waitrequest                               (mm_interconnect_0_fifo_q_5_in_waitrequest),                    //                                                .waitrequest
		.fifo_q_5_in_csr_address                               (mm_interconnect_0_fifo_q_5_in_csr_address),                    //                                 fifo_q_5_in_csr.address
		.fifo_q_5_in_csr_write                                 (mm_interconnect_0_fifo_q_5_in_csr_write),                      //                                                .write
		.fifo_q_5_in_csr_read                                  (mm_interconnect_0_fifo_q_5_in_csr_read),                       //                                                .read
		.fifo_q_5_in_csr_readdata                              (mm_interconnect_0_fifo_q_5_in_csr_readdata),                   //                                                .readdata
		.fifo_q_5_in_csr_writedata                             (mm_interconnect_0_fifo_q_5_in_csr_writedata),                  //                                                .writedata
		.fifo_q_5_out_read                                     (mm_interconnect_0_fifo_q_5_out_read),                          //                                    fifo_q_5_out.read
		.fifo_q_5_out_readdata                                 (mm_interconnect_0_fifo_q_5_out_readdata),                      //                                                .readdata
		.fifo_q_5_out_waitrequest                              (mm_interconnect_0_fifo_q_5_out_waitrequest),                   //                                                .waitrequest
		.fifo_q_6_in_write                                     (mm_interconnect_0_fifo_q_6_in_write),                          //                                     fifo_q_6_in.write
		.fifo_q_6_in_writedata                                 (mm_interconnect_0_fifo_q_6_in_writedata),                      //                                                .writedata
		.fifo_q_6_in_waitrequest                               (mm_interconnect_0_fifo_q_6_in_waitrequest),                    //                                                .waitrequest
		.fifo_q_6_in_csr_address                               (mm_interconnect_0_fifo_q_6_in_csr_address),                    //                                 fifo_q_6_in_csr.address
		.fifo_q_6_in_csr_write                                 (mm_interconnect_0_fifo_q_6_in_csr_write),                      //                                                .write
		.fifo_q_6_in_csr_read                                  (mm_interconnect_0_fifo_q_6_in_csr_read),                       //                                                .read
		.fifo_q_6_in_csr_readdata                              (mm_interconnect_0_fifo_q_6_in_csr_readdata),                   //                                                .readdata
		.fifo_q_6_in_csr_writedata                             (mm_interconnect_0_fifo_q_6_in_csr_writedata),                  //                                                .writedata
		.fifo_q_6_out_read                                     (mm_interconnect_0_fifo_q_6_out_read),                          //                                    fifo_q_6_out.read
		.fifo_q_6_out_readdata                                 (mm_interconnect_0_fifo_q_6_out_readdata),                      //                                                .readdata
		.fifo_q_6_out_waitrequest                              (mm_interconnect_0_fifo_q_6_out_waitrequest),                   //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),        //                     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),          //                                                .write
		.jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),           //                                                .read
		.jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),       //                                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),      //                                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),    //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),     //                                                .chipselect
		.jtag_uart_1b_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_address),     //                  jtag_uart_1b_avalon_jtag_slave.address
		.jtag_uart_1b_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_1b_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_1b_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_1b_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_1b_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_1b_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_1b_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.jtag_uart_1c_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_address),     //                  jtag_uart_1c_avalon_jtag_slave.address
		.jtag_uart_1c_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_1c_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_1c_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_1c_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_1c_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_1c_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_1c_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.jtag_uart_1d_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_address),     //                  jtag_uart_1d_avalon_jtag_slave.address
		.jtag_uart_1d_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_1d_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_1d_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_1d_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_1d_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_1d_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_1d_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.jtag_uart_1e_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_address),     //                  jtag_uart_1e_avalon_jtag_slave.address
		.jtag_uart_1e_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_1e_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_1e_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_1e_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_1e_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_1e_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_1e_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.jtag_uart_1f_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_address),     //                  jtag_uart_1f_avalon_jtag_slave.address
		.jtag_uart_1f_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_1f_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_1f_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_1f_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_1f_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_1f_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.onchip_mem_1b_s1_address                              (mm_interconnect_0_onchip_mem_1b_s1_address),                   //                                onchip_mem_1b_s1.address
		.onchip_mem_1b_s1_write                                (mm_interconnect_0_onchip_mem_1b_s1_write),                     //                                                .write
		.onchip_mem_1b_s1_readdata                             (mm_interconnect_0_onchip_mem_1b_s1_readdata),                  //                                                .readdata
		.onchip_mem_1b_s1_writedata                            (mm_interconnect_0_onchip_mem_1b_s1_writedata),                 //                                                .writedata
		.onchip_mem_1b_s1_byteenable                           (mm_interconnect_0_onchip_mem_1b_s1_byteenable),                //                                                .byteenable
		.onchip_mem_1b_s1_chipselect                           (mm_interconnect_0_onchip_mem_1b_s1_chipselect),                //                                                .chipselect
		.onchip_mem_1b_s1_clken                                (mm_interconnect_0_onchip_mem_1b_s1_clken),                     //                                                .clken
		.onchip_mem_1c_s1_address                              (mm_interconnect_0_onchip_mem_1c_s1_address),                   //                                onchip_mem_1c_s1.address
		.onchip_mem_1c_s1_write                                (mm_interconnect_0_onchip_mem_1c_s1_write),                     //                                                .write
		.onchip_mem_1c_s1_readdata                             (mm_interconnect_0_onchip_mem_1c_s1_readdata),                  //                                                .readdata
		.onchip_mem_1c_s1_writedata                            (mm_interconnect_0_onchip_mem_1c_s1_writedata),                 //                                                .writedata
		.onchip_mem_1c_s1_byteenable                           (mm_interconnect_0_onchip_mem_1c_s1_byteenable),                //                                                .byteenable
		.onchip_mem_1c_s1_chipselect                           (mm_interconnect_0_onchip_mem_1c_s1_chipselect),                //                                                .chipselect
		.onchip_mem_1c_s1_clken                                (mm_interconnect_0_onchip_mem_1c_s1_clken),                     //                                                .clken
		.onchip_mem_1d_s1_address                              (mm_interconnect_0_onchip_mem_1d_s1_address),                   //                                onchip_mem_1d_s1.address
		.onchip_mem_1d_s1_write                                (mm_interconnect_0_onchip_mem_1d_s1_write),                     //                                                .write
		.onchip_mem_1d_s1_readdata                             (mm_interconnect_0_onchip_mem_1d_s1_readdata),                  //                                                .readdata
		.onchip_mem_1d_s1_writedata                            (mm_interconnect_0_onchip_mem_1d_s1_writedata),                 //                                                .writedata
		.onchip_mem_1d_s1_byteenable                           (mm_interconnect_0_onchip_mem_1d_s1_byteenable),                //                                                .byteenable
		.onchip_mem_1d_s1_chipselect                           (mm_interconnect_0_onchip_mem_1d_s1_chipselect),                //                                                .chipselect
		.onchip_mem_1d_s1_clken                                (mm_interconnect_0_onchip_mem_1d_s1_clken),                     //                                                .clken
		.onchip_mem_1e_s1_address                              (mm_interconnect_0_onchip_mem_1e_s1_address),                   //                                onchip_mem_1e_s1.address
		.onchip_mem_1e_s1_write                                (mm_interconnect_0_onchip_mem_1e_s1_write),                     //                                                .write
		.onchip_mem_1e_s1_readdata                             (mm_interconnect_0_onchip_mem_1e_s1_readdata),                  //                                                .readdata
		.onchip_mem_1e_s1_writedata                            (mm_interconnect_0_onchip_mem_1e_s1_writedata),                 //                                                .writedata
		.onchip_mem_1e_s1_byteenable                           (mm_interconnect_0_onchip_mem_1e_s1_byteenable),                //                                                .byteenable
		.onchip_mem_1e_s1_chipselect                           (mm_interconnect_0_onchip_mem_1e_s1_chipselect),                //                                                .chipselect
		.onchip_mem_1e_s1_clken                                (mm_interconnect_0_onchip_mem_1e_s1_clken),                     //                                                .clken
		.onchip_mem_1f_s1_address                              (mm_interconnect_0_onchip_mem_1f_s1_address),                   //                                onchip_mem_1f_s1.address
		.onchip_mem_1f_s1_write                                (mm_interconnect_0_onchip_mem_1f_s1_write),                     //                                                .write
		.onchip_mem_1f_s1_readdata                             (mm_interconnect_0_onchip_mem_1f_s1_readdata),                  //                                                .readdata
		.onchip_mem_1f_s1_writedata                            (mm_interconnect_0_onchip_mem_1f_s1_writedata),                 //                                                .writedata
		.onchip_mem_1f_s1_byteenable                           (mm_interconnect_0_onchip_mem_1f_s1_byteenable),                //                                                .byteenable
		.onchip_mem_1f_s1_chipselect                           (mm_interconnect_0_onchip_mem_1f_s1_chipselect),                //                                                .chipselect
		.onchip_mem_1f_s1_clken                                (mm_interconnect_0_onchip_mem_1f_s1_clken),                     //                                                .clken
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                      //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                        //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                         //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                     //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                    //                                                .writedata
		.sdram_controller_s1_address                           (mm_interconnect_0_sdram_controller_s1_address),                //                             sdram_controller_s1.address
		.sdram_controller_s1_write                             (mm_interconnect_0_sdram_controller_s1_write),                  //                                                .write
		.sdram_controller_s1_read                              (mm_interconnect_0_sdram_controller_s1_read),                   //                                                .read
		.sdram_controller_s1_readdata                          (mm_interconnect_0_sdram_controller_s1_readdata),               //                                                .readdata
		.sdram_controller_s1_writedata                         (mm_interconnect_0_sdram_controller_s1_writedata),              //                                                .writedata
		.sdram_controller_s1_byteenable                        (mm_interconnect_0_sdram_controller_s1_byteenable),             //                                                .byteenable
		.sdram_controller_s1_readdatavalid                     (mm_interconnect_0_sdram_controller_s1_readdatavalid),          //                                                .readdatavalid
		.sdram_controller_s1_waitrequest                       (mm_interconnect_0_sdram_controller_s1_waitrequest),            //                                                .waitrequest
		.sdram_controller_s1_chipselect                        (mm_interconnect_0_sdram_controller_s1_chipselect),             //                                                .chipselect
		.sys_id_control_slave_address                          (mm_interconnect_0_sys_id_control_slave_address),               //                            sys_id_control_slave.address
		.sys_id_control_slave_readdata                         (mm_interconnect_0_sys_id_control_slave_readdata),              //                                                .readdata
		.sysid_1b_control_slave_address                        (mm_interconnect_0_sysid_1b_control_slave_address),             //                          sysid_1b_control_slave.address
		.sysid_1b_control_slave_readdata                       (mm_interconnect_0_sysid_1b_control_slave_readdata),            //                                                .readdata
		.sysid_1c_control_slave_address                        (mm_interconnect_0_sysid_1c_control_slave_address),             //                          sysid_1c_control_slave.address
		.sysid_1c_control_slave_readdata                       (mm_interconnect_0_sysid_1c_control_slave_readdata),            //                                                .readdata
		.sysid_1d_control_slave_address                        (mm_interconnect_0_sysid_1d_control_slave_address),             //                          sysid_1d_control_slave.address
		.sysid_1d_control_slave_readdata                       (mm_interconnect_0_sysid_1d_control_slave_readdata),            //                                                .readdata
		.sysid_1e_control_slave_address                        (mm_interconnect_0_sysid_1e_control_slave_address),             //                          sysid_1e_control_slave.address
		.sysid_1e_control_slave_readdata                       (mm_interconnect_0_sysid_1e_control_slave_readdata),            //                                                .readdata
		.sysid_1f_control_slave_address                        (mm_interconnect_0_sysid_1f_control_slave_address),             //                          sysid_1f_control_slave.address
		.sysid_1f_control_slave_readdata                       (mm_interconnect_0_sysid_1f_control_slave_readdata),            //                                                .readdata
		.timer_s1_address                                      (mm_interconnect_0_timer_s1_address),                           //                                        timer_s1.address
		.timer_s1_write                                        (mm_interconnect_0_timer_s1_write),                             //                                                .write
		.timer_s1_readdata                                     (mm_interconnect_0_timer_s1_readdata),                          //                                                .readdata
		.timer_s1_writedata                                    (mm_interconnect_0_timer_s1_writedata),                         //                                                .writedata
		.timer_s1_chipselect                                   (mm_interconnect_0_timer_s1_chipselect),                        //                                                .chipselect
		.timer_1b_s1_address                                   (mm_interconnect_0_timer_1b_s1_address),                        //                                     timer_1b_s1.address
		.timer_1b_s1_write                                     (mm_interconnect_0_timer_1b_s1_write),                          //                                                .write
		.timer_1b_s1_readdata                                  (mm_interconnect_0_timer_1b_s1_readdata),                       //                                                .readdata
		.timer_1b_s1_writedata                                 (mm_interconnect_0_timer_1b_s1_writedata),                      //                                                .writedata
		.timer_1b_s1_chipselect                                (mm_interconnect_0_timer_1b_s1_chipselect),                     //                                                .chipselect
		.timer_1c_s1_address                                   (mm_interconnect_0_timer_1c_s1_address),                        //                                     timer_1c_s1.address
		.timer_1c_s1_write                                     (mm_interconnect_0_timer_1c_s1_write),                          //                                                .write
		.timer_1c_s1_readdata                                  (mm_interconnect_0_timer_1c_s1_readdata),                       //                                                .readdata
		.timer_1c_s1_writedata                                 (mm_interconnect_0_timer_1c_s1_writedata),                      //                                                .writedata
		.timer_1c_s1_chipselect                                (mm_interconnect_0_timer_1c_s1_chipselect),                     //                                                .chipselect
		.timer_1d_s1_address                                   (mm_interconnect_0_timer_1d_s1_address),                        //                                     timer_1d_s1.address
		.timer_1d_s1_write                                     (mm_interconnect_0_timer_1d_s1_write),                          //                                                .write
		.timer_1d_s1_readdata                                  (mm_interconnect_0_timer_1d_s1_readdata),                       //                                                .readdata
		.timer_1d_s1_writedata                                 (mm_interconnect_0_timer_1d_s1_writedata),                      //                                                .writedata
		.timer_1d_s1_chipselect                                (mm_interconnect_0_timer_1d_s1_chipselect),                     //                                                .chipselect
		.timer_1e_s1_address                                   (mm_interconnect_0_timer_1e_s1_address),                        //                                     timer_1e_s1.address
		.timer_1e_s1_write                                     (mm_interconnect_0_timer_1e_s1_write),                          //                                                .write
		.timer_1e_s1_readdata                                  (mm_interconnect_0_timer_1e_s1_readdata),                       //                                                .readdata
		.timer_1e_s1_writedata                                 (mm_interconnect_0_timer_1e_s1_writedata),                      //                                                .writedata
		.timer_1e_s1_chipselect                                (mm_interconnect_0_timer_1e_s1_chipselect),                     //                                                .chipselect
		.timer_1f_s1_address                                   (mm_interconnect_0_timer_1f_s1_address),                        //                                     timer_1f_s1.address
		.timer_1f_s1_write                                     (mm_interconnect_0_timer_1f_s1_write),                          //                                                .write
		.timer_1f_s1_readdata                                  (mm_interconnect_0_timer_1f_s1_readdata),                       //                                                .readdata
		.timer_1f_s1_writedata                                 (mm_interconnect_0_timer_1f_s1_writedata),                      //                                                .writedata
		.timer_1f_s1_chipselect                                (mm_interconnect_0_timer_1f_s1_chipselect)                      //                                                .chipselect
	);

	Mega_JSoC_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	Mega_JSoC_irq_mapper irq_mapper_001 (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_1b_d_irq_irq)                //    sender.irq
	);

	Mega_JSoC_irq_mapper irq_mapper_002 (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_002_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_1c_d_irq_irq)                //    sender.irq
	);

	Mega_JSoC_irq_mapper irq_mapper_003 (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_003_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_003_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_1d_d_irq_irq)                //    sender.irq
	);

	Mega_JSoC_irq_mapper irq_mapper_004 (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_004_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_004_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_1e_d_irq_irq)                //    sender.irq
	);

	Mega_JSoC_irq_mapper irq_mapper_005 (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_005_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_005_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_1f_d_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (7),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),    // reset_in1.reset
		.reset_in2      (cpu_1b_jtag_debug_module_reset_reset), // reset_in2.reset
		.reset_in3      (cpu_1c_jtag_debug_module_reset_reset), // reset_in3.reset
		.reset_in4      (cpu_1d_jtag_debug_module_reset_reset), // reset_in4.reset
		.reset_in5      (cpu_1e_jtag_debug_module_reset_reset), // reset_in5.reset
		.reset_in6      (cpu_1f_jtag_debug_module_reset_reset), // reset_in6.reset
		.clk            (pll_c0_clk),                           //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (7),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),    // reset_in1.reset
		.reset_in2      (cpu_1b_jtag_debug_module_reset_reset), // reset_in2.reset
		.reset_in3      (cpu_1c_jtag_debug_module_reset_reset), // reset_in3.reset
		.reset_in4      (cpu_1d_jtag_debug_module_reset_reset), // reset_in4.reset
		.reset_in5      (cpu_1e_jtag_debug_module_reset_reset), // reset_in5.reset
		.reset_in6      (cpu_1f_jtag_debug_module_reset_reset), // reset_in6.reset
		.clk            (clk_clk),                              //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

endmodule
