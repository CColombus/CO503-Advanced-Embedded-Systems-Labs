// mpsoc.v

// Generated using ACDS version 13.1 162 at 2024.05.12.18:04:37

`timescale 1 ps / 1 ps
module mpsoc (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire   [0:0] mm_interconnect_0_sysid_1_control_slave_address;             // mm_interconnect_0:sysid_1_control_slave_address -> sysid_1:address
	wire  [31:0] mm_interconnect_0_sysid_1_control_slave_readdata;            // sysid_1:readdata -> mm_interconnect_0:sysid_1_control_slave_readdata
	wire  [31:0] mm_interconnect_0_data_mem_shared_s1_writedata;              // mm_interconnect_0:data_mem_shared_s1_writedata -> data_mem_shared:writedata
	wire  [14:0] mm_interconnect_0_data_mem_shared_s1_address;                // mm_interconnect_0:data_mem_shared_s1_address -> data_mem_shared:address
	wire         mm_interconnect_0_data_mem_shared_s1_chipselect;             // mm_interconnect_0:data_mem_shared_s1_chipselect -> data_mem_shared:chipselect
	wire         mm_interconnect_0_data_mem_shared_s1_clken;                  // mm_interconnect_0:data_mem_shared_s1_clken -> data_mem_shared:clken
	wire         mm_interconnect_0_data_mem_shared_s1_write;                  // mm_interconnect_0:data_mem_shared_s1_write -> data_mem_shared:write
	wire  [31:0] mm_interconnect_0_data_mem_shared_s1_readdata;               // data_mem_shared:readdata -> mm_interconnect_0:data_mem_shared_s1_readdata
	wire   [3:0] mm_interconnect_0_data_mem_shared_s1_byteenable;             // mm_interconnect_0:data_mem_shared_s1_byteenable -> data_mem_shared:byteenable
	wire         mm_interconnect_0_cpu0_jtag_debug_module_waitrequest;        // cpu0:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu0_jtag_debug_module_writedata;          // mm_interconnect_0:cpu0_jtag_debug_module_writedata -> cpu0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu0_jtag_debug_module_address;            // mm_interconnect_0:cpu0_jtag_debug_module_address -> cpu0:jtag_debug_module_address
	wire         mm_interconnect_0_cpu0_jtag_debug_module_write;              // mm_interconnect_0:cpu0_jtag_debug_module_write -> cpu0:jtag_debug_module_write
	wire         mm_interconnect_0_cpu0_jtag_debug_module_read;               // mm_interconnect_0:cpu0_jtag_debug_module_read -> cpu0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu0_jtag_debug_module_readdata;           // cpu0:jtag_debug_module_readdata -> mm_interconnect_0:cpu0_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu0_jtag_debug_module_debugaccess;        // mm_interconnect_0:cpu0_jtag_debug_module_debugaccess -> cpu0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu0_jtag_debug_module_byteenable;         // mm_interconnect_0:cpu0_jtag_debug_module_byteenable -> cpu0:jtag_debug_module_byteenable
	wire         cpu1_instruction_master_waitrequest;                         // mm_interconnect_0:cpu1_instruction_master_waitrequest -> cpu1:i_waitrequest
	wire  [18:0] cpu1_instruction_master_address;                             // cpu1:i_address -> mm_interconnect_0:cpu1_instruction_master_address
	wire         cpu1_instruction_master_read;                                // cpu1:i_read -> mm_interconnect_0:cpu1_instruction_master_read
	wire  [31:0] cpu1_instruction_master_readdata;                            // mm_interconnect_0:cpu1_instruction_master_readdata -> cpu1:i_readdata
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest; // jtag_uart_1:av_waitrequest -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_writedata -> jtag_uart_1:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_address -> jtag_uart_1:av_address
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_chipselect -> jtag_uart_1:av_chipselect
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_write -> jtag_uart_1:av_write_n
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_read -> jtag_uart_1:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata;    // jtag_uart_1:av_readdata -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_ins_mem_c0_s1_writedata;                   // mm_interconnect_0:ins_mem_c0_s1_writedata -> ins_mem_c0:writedata
	wire  [14:0] mm_interconnect_0_ins_mem_c0_s1_address;                     // mm_interconnect_0:ins_mem_c0_s1_address -> ins_mem_c0:address
	wire         mm_interconnect_0_ins_mem_c0_s1_chipselect;                  // mm_interconnect_0:ins_mem_c0_s1_chipselect -> ins_mem_c0:chipselect
	wire         mm_interconnect_0_ins_mem_c0_s1_clken;                       // mm_interconnect_0:ins_mem_c0_s1_clken -> ins_mem_c0:clken
	wire         mm_interconnect_0_ins_mem_c0_s1_write;                       // mm_interconnect_0:ins_mem_c0_s1_write -> ins_mem_c0:write
	wire  [31:0] mm_interconnect_0_ins_mem_c0_s1_readdata;                    // ins_mem_c0:readdata -> mm_interconnect_0:ins_mem_c0_s1_readdata
	wire   [3:0] mm_interconnect_0_ins_mem_c0_s1_byteenable;                  // mm_interconnect_0:ins_mem_c0_s1_byteenable -> ins_mem_c0:byteenable
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire  [31:0] mm_interconnect_0_ins_mem_c1_s1_writedata;                   // mm_interconnect_0:ins_mem_c1_s1_writedata -> ins_mem_c1:writedata
	wire  [14:0] mm_interconnect_0_ins_mem_c1_s1_address;                     // mm_interconnect_0:ins_mem_c1_s1_address -> ins_mem_c1:address
	wire         mm_interconnect_0_ins_mem_c1_s1_chipselect;                  // mm_interconnect_0:ins_mem_c1_s1_chipselect -> ins_mem_c1:chipselect
	wire         mm_interconnect_0_ins_mem_c1_s1_clken;                       // mm_interconnect_0:ins_mem_c1_s1_clken -> ins_mem_c1:clken
	wire         mm_interconnect_0_ins_mem_c1_s1_write;                       // mm_interconnect_0:ins_mem_c1_s1_write -> ins_mem_c1:write
	wire  [31:0] mm_interconnect_0_ins_mem_c1_s1_readdata;                    // ins_mem_c1:readdata -> mm_interconnect_0:ins_mem_c1_s1_readdata
	wire   [3:0] mm_interconnect_0_ins_mem_c1_s1_byteenable;                  // mm_interconnect_0:ins_mem_c1_s1_byteenable -> ins_mem_c1:byteenable
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         cpu0_data_master_waitrequest;                                // mm_interconnect_0:cpu0_data_master_waitrequest -> cpu0:d_waitrequest
	wire  [31:0] cpu0_data_master_writedata;                                  // cpu0:d_writedata -> mm_interconnect_0:cpu0_data_master_writedata
	wire  [19:0] cpu0_data_master_address;                                    // cpu0:d_address -> mm_interconnect_0:cpu0_data_master_address
	wire         cpu0_data_master_write;                                      // cpu0:d_write -> mm_interconnect_0:cpu0_data_master_write
	wire         cpu0_data_master_read;                                       // cpu0:d_read -> mm_interconnect_0:cpu0_data_master_read
	wire  [31:0] cpu0_data_master_readdata;                                   // mm_interconnect_0:cpu0_data_master_readdata -> cpu0:d_readdata
	wire         cpu0_data_master_debugaccess;                                // cpu0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu0_data_master_debugaccess
	wire   [3:0] cpu0_data_master_byteenable;                                 // cpu0:d_byteenable -> mm_interconnect_0:cpu0_data_master_byteenable
	wire         cpu0_instruction_master_waitrequest;                         // mm_interconnect_0:cpu0_instruction_master_waitrequest -> cpu0:i_waitrequest
	wire  [19:0] cpu0_instruction_master_address;                             // cpu0:i_address -> mm_interconnect_0:cpu0_instruction_master_address
	wire         cpu0_instruction_master_read;                                // cpu0:i_read -> mm_interconnect_0:cpu0_instruction_master_read
	wire  [31:0] cpu0_instruction_master_readdata;                            // mm_interconnect_0:cpu0_instruction_master_readdata -> cpu0:i_readdata
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                      // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                        // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_chipselect;                     // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire         mm_interconnect_0_timer_1_s1_write;                          // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                       // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire         mm_interconnect_0_cpu1_jtag_debug_module_waitrequest;        // cpu1:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu1_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu1_jtag_debug_module_writedata;          // mm_interconnect_0:cpu1_jtag_debug_module_writedata -> cpu1:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu1_jtag_debug_module_address;            // mm_interconnect_0:cpu1_jtag_debug_module_address -> cpu1:jtag_debug_module_address
	wire         mm_interconnect_0_cpu1_jtag_debug_module_write;              // mm_interconnect_0:cpu1_jtag_debug_module_write -> cpu1:jtag_debug_module_write
	wire         mm_interconnect_0_cpu1_jtag_debug_module_read;               // mm_interconnect_0:cpu1_jtag_debug_module_read -> cpu1:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu1_jtag_debug_module_readdata;           // cpu1:jtag_debug_module_readdata -> mm_interconnect_0:cpu1_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu1_jtag_debug_module_debugaccess;        // mm_interconnect_0:cpu1_jtag_debug_module_debugaccess -> cpu1:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu1_jtag_debug_module_byteenable;         // mm_interconnect_0:cpu1_jtag_debug_module_byteenable -> cpu1:jtag_debug_module_byteenable
	wire   [0:0] mm_interconnect_0_sysid_0_control_slave_address;             // mm_interconnect_0:sysid_0_control_slave_address -> sysid_0:address
	wire  [31:0] mm_interconnect_0_sysid_0_control_slave_readdata;            // sysid_0:readdata -> mm_interconnect_0:sysid_0_control_slave_readdata
	wire         cpu1_data_master_waitrequest;                                // mm_interconnect_0:cpu1_data_master_waitrequest -> cpu1:d_waitrequest
	wire  [31:0] cpu1_data_master_writedata;                                  // cpu1:d_writedata -> mm_interconnect_0:cpu1_data_master_writedata
	wire  [18:0] cpu1_data_master_address;                                    // cpu1:d_address -> mm_interconnect_0:cpu1_data_master_address
	wire         cpu1_data_master_write;                                      // cpu1:d_write -> mm_interconnect_0:cpu1_data_master_write
	wire         cpu1_data_master_read;                                       // cpu1:d_read -> mm_interconnect_0:cpu1_data_master_read
	wire  [31:0] cpu1_data_master_readdata;                                   // mm_interconnect_0:cpu1_data_master_readdata -> cpu1:d_readdata
	wire         cpu1_data_master_debugaccess;                                // cpu1:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu1_data_master_debugaccess
	wire   [3:0] cpu1_data_master_byteenable;                                 // cpu1:d_byteenable -> mm_interconnect_0:cpu1_data_master_byteenable
	wire         irq_mapper_receiver0_irq;                                    // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu0_d_irq_irq;                                              // irq_mapper:sender_irq -> cpu0:d_irq
	wire         irq_mapper_001_receiver0_irq;                                // timer_1:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                // jtag_uart_1:av_irq -> irq_mapper_001:receiver1_irq
	wire  [31:0] cpu1_d_irq_irq;                                              // irq_mapper_001:sender_irq -> cpu1:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [cpu0:reset_n, ins_mem_c0:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:cpu0_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, sysid_0:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu0:reset_req, ins_mem_c0:reset_req, rst_translator:reset_req_in]
	wire         cpu0_jtag_debug_module_reset_reset;                          // cpu0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in2]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [data_mem_shared:reset, mm_interconnect_0:data_mem_shared_reset1_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> data_mem_shared:reset_req
	wire         cpu1_jtag_debug_module_reset_reset;                          // cpu1:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [cpu1:reset_n, ins_mem_c1:reset, irq_mapper_001:reset, jtag_uart_1:rst_n, mm_interconnect_0:cpu1_reset_n_reset_bridge_in_reset_reset, rst_translator_002:in_reset, sysid_1:reset_n, timer_1:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                      // rst_controller_002:reset_req -> [cpu1:reset_req, ins_mem_c1:reset_req, rst_translator_002:reset_req_in]

	mpsoc_ins_mem_c0 ins_mem_c0 (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_ins_mem_c0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ins_mem_c0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ins_mem_c0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ins_mem_c0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ins_mem_c0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ins_mem_c0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ins_mem_c0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	mpsoc_cpu0 cpu0 (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (cpu0_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu0_data_master_read),                                //                          .read
		.d_readdata                            (cpu0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu0_data_master_write),                               //                          .write
		.d_writedata                           (cpu0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu0_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	mpsoc_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	mpsoc_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	mpsoc_sysid_0 sysid_0 (
		.clock    (clk_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_0_control_slave_address)   //              .address
	);

	mpsoc_data_mem_shared data_mem_shared (
		.clk        (clk_clk),                                         //   clk1.clk
		.address    (mm_interconnect_0_data_mem_shared_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_mem_shared_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_mem_shared_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_mem_shared_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_mem_shared_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_mem_shared_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_mem_shared_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),              // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)           //       .reset_req
	);

	mpsoc_ins_mem_c1 ins_mem_c1 (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_ins_mem_c1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ins_mem_c1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ins_mem_c1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ins_mem_c1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ins_mem_c1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ins_mem_c1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ins_mem_c1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)      //       .reset_req
	);

	mpsoc_cpu1 cpu1 (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                  //                   reset_n.reset_n
		.reset_req                             (rst_controller_002_reset_out_reset_req),               //                          .reset_req
		.d_address                             (cpu1_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu1_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu1_data_master_read),                                //                          .read
		.d_readdata                            (cpu1_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu1_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu1_data_master_write),                               //                          .write
		.d_writedata                           (cpu1_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu1_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu1_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu1_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu1_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu1_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu1_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu1_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu1_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu1_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu1_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu1_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu1_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu1_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu1_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu1_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	mpsoc_jtag_uart_0 jtag_uart_1 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver1_irq)                                 //               irq.irq
	);

	mpsoc_timer_0 timer_1 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver0_irq)             //   irq.irq
	);

	mpsoc_sysid_1 sysid_1 (
		.clock    (clk_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),              //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_1_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_1_control_slave_address)   //              .address
	);

	mpsoc_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                      (clk_clk),                                                     //                                    clock_clk.clk
		.cpu0_reset_n_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                              //           cpu0_reset_n_reset_bridge_in_reset.reset
		.cpu1_reset_n_reset_bridge_in_reset_reset           (rst_controller_002_reset_out_reset),                          //           cpu1_reset_n_reset_bridge_in_reset.reset
		.data_mem_shared_reset1_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // data_mem_shared_reset1_reset_bridge_in_reset.reset
		.cpu0_data_master_address                           (cpu0_data_master_address),                                    //                             cpu0_data_master.address
		.cpu0_data_master_waitrequest                       (cpu0_data_master_waitrequest),                                //                                             .waitrequest
		.cpu0_data_master_byteenable                        (cpu0_data_master_byteenable),                                 //                                             .byteenable
		.cpu0_data_master_read                              (cpu0_data_master_read),                                       //                                             .read
		.cpu0_data_master_readdata                          (cpu0_data_master_readdata),                                   //                                             .readdata
		.cpu0_data_master_write                             (cpu0_data_master_write),                                      //                                             .write
		.cpu0_data_master_writedata                         (cpu0_data_master_writedata),                                  //                                             .writedata
		.cpu0_data_master_debugaccess                       (cpu0_data_master_debugaccess),                                //                                             .debugaccess
		.cpu0_instruction_master_address                    (cpu0_instruction_master_address),                             //                      cpu0_instruction_master.address
		.cpu0_instruction_master_waitrequest                (cpu0_instruction_master_waitrequest),                         //                                             .waitrequest
		.cpu0_instruction_master_read                       (cpu0_instruction_master_read),                                //                                             .read
		.cpu0_instruction_master_readdata                   (cpu0_instruction_master_readdata),                            //                                             .readdata
		.cpu1_data_master_address                           (cpu1_data_master_address),                                    //                             cpu1_data_master.address
		.cpu1_data_master_waitrequest                       (cpu1_data_master_waitrequest),                                //                                             .waitrequest
		.cpu1_data_master_byteenable                        (cpu1_data_master_byteenable),                                 //                                             .byteenable
		.cpu1_data_master_read                              (cpu1_data_master_read),                                       //                                             .read
		.cpu1_data_master_readdata                          (cpu1_data_master_readdata),                                   //                                             .readdata
		.cpu1_data_master_write                             (cpu1_data_master_write),                                      //                                             .write
		.cpu1_data_master_writedata                         (cpu1_data_master_writedata),                                  //                                             .writedata
		.cpu1_data_master_debugaccess                       (cpu1_data_master_debugaccess),                                //                                             .debugaccess
		.cpu1_instruction_master_address                    (cpu1_instruction_master_address),                             //                      cpu1_instruction_master.address
		.cpu1_instruction_master_waitrequest                (cpu1_instruction_master_waitrequest),                         //                                             .waitrequest
		.cpu1_instruction_master_read                       (cpu1_instruction_master_read),                                //                                             .read
		.cpu1_instruction_master_readdata                   (cpu1_instruction_master_readdata),                            //                                             .readdata
		.cpu0_jtag_debug_module_address                     (mm_interconnect_0_cpu0_jtag_debug_module_address),            //                       cpu0_jtag_debug_module.address
		.cpu0_jtag_debug_module_write                       (mm_interconnect_0_cpu0_jtag_debug_module_write),              //                                             .write
		.cpu0_jtag_debug_module_read                        (mm_interconnect_0_cpu0_jtag_debug_module_read),               //                                             .read
		.cpu0_jtag_debug_module_readdata                    (mm_interconnect_0_cpu0_jtag_debug_module_readdata),           //                                             .readdata
		.cpu0_jtag_debug_module_writedata                   (mm_interconnect_0_cpu0_jtag_debug_module_writedata),          //                                             .writedata
		.cpu0_jtag_debug_module_byteenable                  (mm_interconnect_0_cpu0_jtag_debug_module_byteenable),         //                                             .byteenable
		.cpu0_jtag_debug_module_waitrequest                 (mm_interconnect_0_cpu0_jtag_debug_module_waitrequest),        //                                             .waitrequest
		.cpu0_jtag_debug_module_debugaccess                 (mm_interconnect_0_cpu0_jtag_debug_module_debugaccess),        //                                             .debugaccess
		.cpu1_jtag_debug_module_address                     (mm_interconnect_0_cpu1_jtag_debug_module_address),            //                       cpu1_jtag_debug_module.address
		.cpu1_jtag_debug_module_write                       (mm_interconnect_0_cpu1_jtag_debug_module_write),              //                                             .write
		.cpu1_jtag_debug_module_read                        (mm_interconnect_0_cpu1_jtag_debug_module_read),               //                                             .read
		.cpu1_jtag_debug_module_readdata                    (mm_interconnect_0_cpu1_jtag_debug_module_readdata),           //                                             .readdata
		.cpu1_jtag_debug_module_writedata                   (mm_interconnect_0_cpu1_jtag_debug_module_writedata),          //                                             .writedata
		.cpu1_jtag_debug_module_byteenable                  (mm_interconnect_0_cpu1_jtag_debug_module_byteenable),         //                                             .byteenable
		.cpu1_jtag_debug_module_waitrequest                 (mm_interconnect_0_cpu1_jtag_debug_module_waitrequest),        //                                             .waitrequest
		.cpu1_jtag_debug_module_debugaccess                 (mm_interconnect_0_cpu1_jtag_debug_module_debugaccess),        //                                             .debugaccess
		.data_mem_shared_s1_address                         (mm_interconnect_0_data_mem_shared_s1_address),                //                           data_mem_shared_s1.address
		.data_mem_shared_s1_write                           (mm_interconnect_0_data_mem_shared_s1_write),                  //                                             .write
		.data_mem_shared_s1_readdata                        (mm_interconnect_0_data_mem_shared_s1_readdata),               //                                             .readdata
		.data_mem_shared_s1_writedata                       (mm_interconnect_0_data_mem_shared_s1_writedata),              //                                             .writedata
		.data_mem_shared_s1_byteenable                      (mm_interconnect_0_data_mem_shared_s1_byteenable),             //                                             .byteenable
		.data_mem_shared_s1_chipselect                      (mm_interconnect_0_data_mem_shared_s1_chipselect),             //                                             .chipselect
		.data_mem_shared_s1_clken                           (mm_interconnect_0_data_mem_shared_s1_clken),                  //                                             .clken
		.ins_mem_c0_s1_address                              (mm_interconnect_0_ins_mem_c0_s1_address),                     //                                ins_mem_c0_s1.address
		.ins_mem_c0_s1_write                                (mm_interconnect_0_ins_mem_c0_s1_write),                       //                                             .write
		.ins_mem_c0_s1_readdata                             (mm_interconnect_0_ins_mem_c0_s1_readdata),                    //                                             .readdata
		.ins_mem_c0_s1_writedata                            (mm_interconnect_0_ins_mem_c0_s1_writedata),                   //                                             .writedata
		.ins_mem_c0_s1_byteenable                           (mm_interconnect_0_ins_mem_c0_s1_byteenable),                  //                                             .byteenable
		.ins_mem_c0_s1_chipselect                           (mm_interconnect_0_ins_mem_c0_s1_chipselect),                  //                                             .chipselect
		.ins_mem_c0_s1_clken                                (mm_interconnect_0_ins_mem_c0_s1_clken),                       //                                             .clken
		.ins_mem_c1_s1_address                              (mm_interconnect_0_ins_mem_c1_s1_address),                     //                                ins_mem_c1_s1.address
		.ins_mem_c1_s1_write                                (mm_interconnect_0_ins_mem_c1_s1_write),                       //                                             .write
		.ins_mem_c1_s1_readdata                             (mm_interconnect_0_ins_mem_c1_s1_readdata),                    //                                             .readdata
		.ins_mem_c1_s1_writedata                            (mm_interconnect_0_ins_mem_c1_s1_writedata),                   //                                             .writedata
		.ins_mem_c1_s1_byteenable                           (mm_interconnect_0_ins_mem_c1_s1_byteenable),                  //                                             .byteenable
		.ins_mem_c1_s1_chipselect                           (mm_interconnect_0_ins_mem_c1_s1_chipselect),                  //                                             .chipselect
		.ins_mem_c1_s1_clken                                (mm_interconnect_0_ins_mem_c1_s1_clken),                       //                                             .clken
		.jtag_uart_0_avalon_jtag_slave_address              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                             .write
		.jtag_uart_0_avalon_jtag_slave_read                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                             .read
		.jtag_uart_0_avalon_jtag_slave_readdata             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                             .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                             .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                             .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                             .chipselect
		.jtag_uart_1_avalon_jtag_slave_address              (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),     //                jtag_uart_1_avalon_jtag_slave.address
		.jtag_uart_1_avalon_jtag_slave_write                (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),       //                                             .write
		.jtag_uart_1_avalon_jtag_slave_read                 (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),        //                                             .read
		.jtag_uart_1_avalon_jtag_slave_readdata             (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),    //                                             .readdata
		.jtag_uart_1_avalon_jtag_slave_writedata            (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),   //                                             .writedata
		.jtag_uart_1_avalon_jtag_slave_waitrequest          (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest), //                                             .waitrequest
		.jtag_uart_1_avalon_jtag_slave_chipselect           (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),  //                                             .chipselect
		.sysid_0_control_slave_address                      (mm_interconnect_0_sysid_0_control_slave_address),             //                        sysid_0_control_slave.address
		.sysid_0_control_slave_readdata                     (mm_interconnect_0_sysid_0_control_slave_readdata),            //                                             .readdata
		.sysid_1_control_slave_address                      (mm_interconnect_0_sysid_1_control_slave_address),             //                        sysid_1_control_slave.address
		.sysid_1_control_slave_readdata                     (mm_interconnect_0_sysid_1_control_slave_readdata),            //                                             .readdata
		.timer_0_s1_address                                 (mm_interconnect_0_timer_0_s1_address),                        //                                   timer_0_s1.address
		.timer_0_s1_write                                   (mm_interconnect_0_timer_0_s1_write),                          //                                             .write
		.timer_0_s1_readdata                                (mm_interconnect_0_timer_0_s1_readdata),                       //                                             .readdata
		.timer_0_s1_writedata                               (mm_interconnect_0_timer_0_s1_writedata),                      //                                             .writedata
		.timer_0_s1_chipselect                              (mm_interconnect_0_timer_0_s1_chipselect),                     //                                             .chipselect
		.timer_1_s1_address                                 (mm_interconnect_0_timer_1_s1_address),                        //                                   timer_1_s1.address
		.timer_1_s1_write                                   (mm_interconnect_0_timer_1_s1_write),                          //                                             .write
		.timer_1_s1_readdata                                (mm_interconnect_0_timer_1_s1_readdata),                       //                                             .readdata
		.timer_1_s1_writedata                               (mm_interconnect_0_timer_1_s1_writedata),                      //                                             .writedata
		.timer_1_s1_chipselect                              (mm_interconnect_0_timer_1_s1_chipselect)                      //                                             .chipselect
	);

	mpsoc_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu0_d_irq_irq)                  //    sender.irq
	);

	mpsoc_irq_mapper irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu1_d_irq_irq)                      //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu1_jtag_debug_module_reset_reset),     // reset_in1.reset
		.reset_in2      (cpu0_jtag_debug_module_reset_reset),     // reset_in2.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu1_jtag_debug_module_reset_reset),     // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
