// FTOP_MSOC_CPU_1b_p2.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module FTOP_MSOC_CPU_1b_p2 (
		input  wire        clock_bridge_0_in_clk_clk,     //   clock_bridge_0_in_clk.clk
		input  wire        mm_bridge_0_m0_waitrequest,    //          mm_bridge_0_m0.waitrequest
		input  wire [31:0] mm_bridge_0_m0_readdata,       //                        .readdata
		input  wire        mm_bridge_0_m0_readdatavalid,  //                        .readdatavalid
		output wire [0:0]  mm_bridge_0_m0_burstcount,     //                        .burstcount
		output wire [31:0] mm_bridge_0_m0_writedata,      //                        .writedata
		output wire [6:0]  mm_bridge_0_m0_address,        //                        .address
		output wire        mm_bridge_0_m0_write,          //                        .write
		output wire        mm_bridge_0_m0_read,           //                        .read
		output wire [3:0]  mm_bridge_0_m0_byteenable,     //                        .byteenable
		output wire        mm_bridge_0_m0_debugaccess,    //                        .debugaccess
		input  wire        reset_bridge_0_in_reset_reset  // reset_bridge_0_in_reset.reset
	);

	wire  [31:0] sub_cpu_0_data_master_readdata;                          // mm_interconnect_0:sub_cpu_0_data_master_readdata -> sub_cpu_0:d_readdata
	wire         sub_cpu_0_data_master_waitrequest;                       // mm_interconnect_0:sub_cpu_0_data_master_waitrequest -> sub_cpu_0:d_waitrequest
	wire         sub_cpu_0_data_master_debugaccess;                       // sub_cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:sub_cpu_0_data_master_debugaccess
	wire  [28:0] sub_cpu_0_data_master_address;                           // sub_cpu_0:d_address -> mm_interconnect_0:sub_cpu_0_data_master_address
	wire   [3:0] sub_cpu_0_data_master_byteenable;                        // sub_cpu_0:d_byteenable -> mm_interconnect_0:sub_cpu_0_data_master_byteenable
	wire         sub_cpu_0_data_master_read;                              // sub_cpu_0:d_read -> mm_interconnect_0:sub_cpu_0_data_master_read
	wire         sub_cpu_0_data_master_write;                             // sub_cpu_0:d_write -> mm_interconnect_0:sub_cpu_0_data_master_write
	wire  [31:0] sub_cpu_0_data_master_writedata;                         // sub_cpu_0:d_writedata -> mm_interconnect_0:sub_cpu_0_data_master_writedata
	wire  [31:0] sub_cpu_0_instruction_master_readdata;                   // mm_interconnect_0:sub_cpu_0_instruction_master_readdata -> sub_cpu_0:i_readdata
	wire         sub_cpu_0_instruction_master_waitrequest;                // mm_interconnect_0:sub_cpu_0_instruction_master_waitrequest -> sub_cpu_0:i_waitrequest
	wire  [16:0] sub_cpu_0_instruction_master_address;                    // sub_cpu_0:i_address -> mm_interconnect_0:sub_cpu_0_instruction_master_address
	wire         sub_cpu_0_instruction_master_read;                       // sub_cpu_0:i_read -> mm_interconnect_0:sub_cpu_0_instruction_master_read
	wire         mm_interconnect_0_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:uart_0_avalon_jtag_slave_chipselect -> uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_uart_0_avalon_jtag_slave_readdata;     // uart_0:av_readdata -> mm_interconnect_0:uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_uart_0_avalon_jtag_slave_waitrequest;  // uart_0:av_waitrequest -> mm_interconnect_0:uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:uart_0_avalon_jtag_slave_address -> uart_0:av_address
	wire         mm_interconnect_0_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:uart_0_avalon_jtag_slave_read -> uart_0:av_read_n
	wire         mm_interconnect_0_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:uart_0_avalon_jtag_slave_write -> uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:uart_0_avalon_jtag_slave_writedata -> uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sub_cpu_0_debug_mem_slave_readdata;    // sub_cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:sub_cpu_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_sub_cpu_0_debug_mem_slave_waitrequest; // sub_cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:sub_cpu_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_sub_cpu_0_debug_mem_slave_debugaccess; // mm_interconnect_0:sub_cpu_0_debug_mem_slave_debugaccess -> sub_cpu_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_sub_cpu_0_debug_mem_slave_address;     // mm_interconnect_0:sub_cpu_0_debug_mem_slave_address -> sub_cpu_0:debug_mem_slave_address
	wire         mm_interconnect_0_sub_cpu_0_debug_mem_slave_read;        // mm_interconnect_0:sub_cpu_0_debug_mem_slave_read -> sub_cpu_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_sub_cpu_0_debug_mem_slave_byteenable;  // mm_interconnect_0:sub_cpu_0_debug_mem_slave_byteenable -> sub_cpu_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_sub_cpu_0_debug_mem_slave_write;       // mm_interconnect_0:sub_cpu_0_debug_mem_slave_write -> sub_cpu_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_sub_cpu_0_debug_mem_slave_writedata;   // mm_interconnect_0:sub_cpu_0_debug_mem_slave_writedata -> sub_cpu_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_readdata;               // mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_bridge_0_s0_waitrequest;            // mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	wire         mm_interconnect_0_mm_bridge_0_s0_debugaccess;            // mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire   [6:0] mm_interconnect_0_mm_bridge_0_s0_address;                // mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_0_mm_bridge_0_s0_read;                   // mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire   [3:0] mm_interconnect_0_mm_bridge_0_s0_byteenable;             // mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire         mm_interconnect_0_mm_bridge_0_s0_readdatavalid;          // mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	wire         mm_interconnect_0_mm_bridge_0_s0_write;                  // mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_writedata;              // mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_bridge_0_s0_burstcount;             // mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire         mm_interconnect_0_oc_ram_0_s1_chipselect;                // mm_interconnect_0:oc_ram_0_s1_chipselect -> oc_ram_0:chipselect
	wire  [31:0] mm_interconnect_0_oc_ram_0_s1_readdata;                  // oc_ram_0:readdata -> mm_interconnect_0:oc_ram_0_s1_readdata
	wire  [12:0] mm_interconnect_0_oc_ram_0_s1_address;                   // mm_interconnect_0:oc_ram_0_s1_address -> oc_ram_0:address
	wire   [3:0] mm_interconnect_0_oc_ram_0_s1_byteenable;                // mm_interconnect_0:oc_ram_0_s1_byteenable -> oc_ram_0:byteenable
	wire         mm_interconnect_0_oc_ram_0_s1_write;                     // mm_interconnect_0:oc_ram_0_s1_write -> oc_ram_0:write
	wire  [31:0] mm_interconnect_0_oc_ram_0_s1_writedata;                 // mm_interconnect_0:oc_ram_0_s1_writedata -> oc_ram_0:writedata
	wire         mm_interconnect_0_oc_ram_0_s1_clken;                     // mm_interconnect_0:oc_ram_0_s1_clken -> oc_ram_0:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                 // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                   // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                    // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                      // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                  // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver0_irq;                                // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                // uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] sub_cpu_0_irq_irq;                                       // irq_mapper:sender_irq -> sub_cpu_0:irq
	wire         rst_controller_reset_out_reset;                          // rst_controller:reset_out -> [irq_mapper:reset, mm_bridge_0:reset, mm_interconnect_0:sub_cpu_0_reset_reset_bridge_in_reset_reset, oc_ram_0:reset, rst_translator:in_reset, sub_cpu_0:reset_n, timer_0:reset_n, uart_0:rst_n]
	wire         rst_controller_reset_out_reset_req;                      // rst_controller:reset_req -> [oc_ram_0:reset_req, rst_translator:reset_req_in, sub_cpu_0:reset_req]
	wire         sub_cpu_0_debug_reset_request_reset;                     // sub_cpu_0:debug_reset_request -> rst_controller:reset_in0

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (7),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clock_bridge_0_in_clk_clk),                      //   clk.clk
		.reset            (rst_controller_reset_out_reset),                 // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	FTOP_MSOC_CPU_1b_p2_oc_ram_0 oc_ram_0 (
		.clk        (clock_bridge_0_in_clk_clk),                //   clk1.clk
		.address    (mm_interconnect_0_oc_ram_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_oc_ram_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_oc_ram_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_oc_ram_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_oc_ram_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_oc_ram_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_oc_ram_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze     (1'b0)                                      // (terminated)
	);

	FTOP_MSOC_CPU_1b_p2_sub_cpu_0 sub_cpu_0 (
		.clk                                 (clock_bridge_0_in_clk_clk),                               //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                         //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                           (sub_cpu_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (sub_cpu_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (sub_cpu_0_data_master_read),                              //                          .read
		.d_readdata                          (sub_cpu_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (sub_cpu_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (sub_cpu_0_data_master_write),                             //                          .write
		.d_writedata                         (sub_cpu_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (sub_cpu_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (sub_cpu_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (sub_cpu_0_instruction_master_read),                       //                          .read
		.i_readdata                          (sub_cpu_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (sub_cpu_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (sub_cpu_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (sub_cpu_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_sub_cpu_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_sub_cpu_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_sub_cpu_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_sub_cpu_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_sub_cpu_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_sub_cpu_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_sub_cpu_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_sub_cpu_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	FTOP_MSOC_timer_1a timer_0 (
		.clk        (clock_bridge_0_in_clk_clk),               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	FTOP_MSOC_jtag_uart_1a uart_0 (
		.clk            (clock_bridge_0_in_clk_clk),                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                        //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                //               irq.irq
	);

	FTOP_MSOC_CPU_1b_p2_mm_interconnect_0 mm_interconnect_0 (
		.clock_bridge_0_out_clk_clk                  (clock_bridge_0_in_clk_clk),                               //                clock_bridge_0_out_clk.clk
		.sub_cpu_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                          // sub_cpu_0_reset_reset_bridge_in_reset.reset
		.sub_cpu_0_data_master_address               (sub_cpu_0_data_master_address),                           //                 sub_cpu_0_data_master.address
		.sub_cpu_0_data_master_waitrequest           (sub_cpu_0_data_master_waitrequest),                       //                                      .waitrequest
		.sub_cpu_0_data_master_byteenable            (sub_cpu_0_data_master_byteenable),                        //                                      .byteenable
		.sub_cpu_0_data_master_read                  (sub_cpu_0_data_master_read),                              //                                      .read
		.sub_cpu_0_data_master_readdata              (sub_cpu_0_data_master_readdata),                          //                                      .readdata
		.sub_cpu_0_data_master_write                 (sub_cpu_0_data_master_write),                             //                                      .write
		.sub_cpu_0_data_master_writedata             (sub_cpu_0_data_master_writedata),                         //                                      .writedata
		.sub_cpu_0_data_master_debugaccess           (sub_cpu_0_data_master_debugaccess),                       //                                      .debugaccess
		.sub_cpu_0_instruction_master_address        (sub_cpu_0_instruction_master_address),                    //          sub_cpu_0_instruction_master.address
		.sub_cpu_0_instruction_master_waitrequest    (sub_cpu_0_instruction_master_waitrequest),                //                                      .waitrequest
		.sub_cpu_0_instruction_master_read           (sub_cpu_0_instruction_master_read),                       //                                      .read
		.sub_cpu_0_instruction_master_readdata       (sub_cpu_0_instruction_master_readdata),                   //                                      .readdata
		.mm_bridge_0_s0_address                      (mm_interconnect_0_mm_bridge_0_s0_address),                //                        mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                        (mm_interconnect_0_mm_bridge_0_s0_write),                  //                                      .write
		.mm_bridge_0_s0_read                         (mm_interconnect_0_mm_bridge_0_s0_read),                   //                                      .read
		.mm_bridge_0_s0_readdata                     (mm_interconnect_0_mm_bridge_0_s0_readdata),               //                                      .readdata
		.mm_bridge_0_s0_writedata                    (mm_interconnect_0_mm_bridge_0_s0_writedata),              //                                      .writedata
		.mm_bridge_0_s0_burstcount                   (mm_interconnect_0_mm_bridge_0_s0_burstcount),             //                                      .burstcount
		.mm_bridge_0_s0_byteenable                   (mm_interconnect_0_mm_bridge_0_s0_byteenable),             //                                      .byteenable
		.mm_bridge_0_s0_readdatavalid                (mm_interconnect_0_mm_bridge_0_s0_readdatavalid),          //                                      .readdatavalid
		.mm_bridge_0_s0_waitrequest                  (mm_interconnect_0_mm_bridge_0_s0_waitrequest),            //                                      .waitrequest
		.mm_bridge_0_s0_debugaccess                  (mm_interconnect_0_mm_bridge_0_s0_debugaccess),            //                                      .debugaccess
		.oc_ram_0_s1_address                         (mm_interconnect_0_oc_ram_0_s1_address),                   //                           oc_ram_0_s1.address
		.oc_ram_0_s1_write                           (mm_interconnect_0_oc_ram_0_s1_write),                     //                                      .write
		.oc_ram_0_s1_readdata                        (mm_interconnect_0_oc_ram_0_s1_readdata),                  //                                      .readdata
		.oc_ram_0_s1_writedata                       (mm_interconnect_0_oc_ram_0_s1_writedata),                 //                                      .writedata
		.oc_ram_0_s1_byteenable                      (mm_interconnect_0_oc_ram_0_s1_byteenable),                //                                      .byteenable
		.oc_ram_0_s1_chipselect                      (mm_interconnect_0_oc_ram_0_s1_chipselect),                //                                      .chipselect
		.oc_ram_0_s1_clken                           (mm_interconnect_0_oc_ram_0_s1_clken),                     //                                      .clken
		.sub_cpu_0_debug_mem_slave_address           (mm_interconnect_0_sub_cpu_0_debug_mem_slave_address),     //             sub_cpu_0_debug_mem_slave.address
		.sub_cpu_0_debug_mem_slave_write             (mm_interconnect_0_sub_cpu_0_debug_mem_slave_write),       //                                      .write
		.sub_cpu_0_debug_mem_slave_read              (mm_interconnect_0_sub_cpu_0_debug_mem_slave_read),        //                                      .read
		.sub_cpu_0_debug_mem_slave_readdata          (mm_interconnect_0_sub_cpu_0_debug_mem_slave_readdata),    //                                      .readdata
		.sub_cpu_0_debug_mem_slave_writedata         (mm_interconnect_0_sub_cpu_0_debug_mem_slave_writedata),   //                                      .writedata
		.sub_cpu_0_debug_mem_slave_byteenable        (mm_interconnect_0_sub_cpu_0_debug_mem_slave_byteenable),  //                                      .byteenable
		.sub_cpu_0_debug_mem_slave_waitrequest       (mm_interconnect_0_sub_cpu_0_debug_mem_slave_waitrequest), //                                      .waitrequest
		.sub_cpu_0_debug_mem_slave_debugaccess       (mm_interconnect_0_sub_cpu_0_debug_mem_slave_debugaccess), //                                      .debugaccess
		.timer_0_s1_address                          (mm_interconnect_0_timer_0_s1_address),                    //                            timer_0_s1.address
		.timer_0_s1_write                            (mm_interconnect_0_timer_0_s1_write),                      //                                      .write
		.timer_0_s1_readdata                         (mm_interconnect_0_timer_0_s1_readdata),                   //                                      .readdata
		.timer_0_s1_writedata                        (mm_interconnect_0_timer_0_s1_writedata),                  //                                      .writedata
		.timer_0_s1_chipselect                       (mm_interconnect_0_timer_0_s1_chipselect),                 //                                      .chipselect
		.uart_0_avalon_jtag_slave_address            (mm_interconnect_0_uart_0_avalon_jtag_slave_address),      //              uart_0_avalon_jtag_slave.address
		.uart_0_avalon_jtag_slave_write              (mm_interconnect_0_uart_0_avalon_jtag_slave_write),        //                                      .write
		.uart_0_avalon_jtag_slave_read               (mm_interconnect_0_uart_0_avalon_jtag_slave_read),         //                                      .read
		.uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_uart_0_avalon_jtag_slave_readdata),     //                                      .readdata
		.uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_uart_0_avalon_jtag_slave_writedata),    //                                      .writedata
		.uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_uart_0_avalon_jtag_slave_waitrequest),  //                                      .waitrequest
		.uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_uart_0_avalon_jtag_slave_chipselect)    //                                      .chipselect
	);

	FTOP_MSOC_irq_mapper irq_mapper (
		.clk           (clock_bridge_0_in_clk_clk),      //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (sub_cpu_0_irq_irq)               //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (sub_cpu_0_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (reset_bridge_0_in_reset_reset),       // reset_in1.reset
		.clk            (clock_bridge_0_in_clk_clk),           //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
