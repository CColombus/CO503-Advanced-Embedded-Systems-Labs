// FTOP_MSOC.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module FTOP_MSOC (
		input  wire        clk_clk,                     //                   clk.clk
		input  wire        reset_reset_n,               //                 reset.reset_n
		output wire        sdram_clk_clk,               //             sdram_clk.clk
		output wire [12:0] sdram_controller_wire_addr,  // sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,    //                      .ba
		output wire        sdram_controller_wire_cas_n, //                      .cas_n
		output wire        sdram_controller_wire_cke,   //                      .cke
		output wire        sdram_controller_wire_cs_n,  //                      .cs_n
		inout  wire [31:0] sdram_controller_wire_dq,    //                      .dq
		output wire [3:0]  sdram_controller_wire_dqm,   //                      .dqm
		output wire        sdram_controller_wire_ras_n, //                      .ras_n
		output wire        sdram_controller_wire_we_n   //                      .we_n
	);

	wire         pll_c0_clk;                                                   // pll:c0 -> [CPU_1b_p1:clock_bridge_0_in_clk_clk, CPU_1b_p2:clock_bridge_0_in_clk_clk, CPU_1b_p3:clock_bridge_0_in_clk_clk, CPU_1c_p1:clock_bridge_0_in_clk_clk, CPU_1c_p2:clock_bridge_0_in_clk_clk, CPU_1c_p3:clock_bridge_0_in_clk_clk, CPU_1d_p1:clock_bridge_0_in_clk_clk, CPU_1d_p2:clock_bridge_0_in_clk_clk, CPU_1d_p3:clock_bridge_0_in_clk_clk, CPU_1e:clock_bridge_0_in_clk_clk, cpu_1a:clk, cpu_1f:clk, fifo_qa_p1:wrclock, fifo_qa_p2:wrclock, fifo_qa_p3:wrclock, fifo_qb_p1:wrclock, fifo_qb_p2:wrclock, fifo_qb_p3:wrclock, fifo_qc_p1:wrclock, fifo_qc_p2:wrclock, fifo_qc_p3:wrclock, fifo_qd_p1:wrclock, fifo_qd_p2:wrclock, fifo_qd_p3:wrclock, fifo_qe:wrclock, irq_mapper:clk, irq_mapper_001:clk, jtag_uart_1a:clk, jtag_uart_1f:clk, mem_info:clk, mm_interconnect_0:pll_c0_clk, oc_ram_1f:clk, rst_controller:clk, sdram_controller:clk, sys_id_1a:clock, sysid_1f:clock, timer_1a:clk, timer_1f:clk]
	wire  [31:0] cpu_1a_data_master_readdata;                                  // mm_interconnect_0:cpu_1a_data_master_readdata -> cpu_1a:d_readdata
	wire         cpu_1a_data_master_waitrequest;                               // mm_interconnect_0:cpu_1a_data_master_waitrequest -> cpu_1a:d_waitrequest
	wire         cpu_1a_data_master_debugaccess;                               // cpu_1a:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1a_data_master_debugaccess
	wire  [27:0] cpu_1a_data_master_address;                                   // cpu_1a:d_address -> mm_interconnect_0:cpu_1a_data_master_address
	wire   [3:0] cpu_1a_data_master_byteenable;                                // cpu_1a:d_byteenable -> mm_interconnect_0:cpu_1a_data_master_byteenable
	wire         cpu_1a_data_master_read;                                      // cpu_1a:d_read -> mm_interconnect_0:cpu_1a_data_master_read
	wire         cpu_1a_data_master_write;                                     // cpu_1a:d_write -> mm_interconnect_0:cpu_1a_data_master_write
	wire  [31:0] cpu_1a_data_master_writedata;                                 // cpu_1a:d_writedata -> mm_interconnect_0:cpu_1a_data_master_writedata
	wire  [31:0] cpu_1f_data_master_readdata;                                  // mm_interconnect_0:cpu_1f_data_master_readdata -> cpu_1f:d_readdata
	wire         cpu_1f_data_master_waitrequest;                               // mm_interconnect_0:cpu_1f_data_master_waitrequest -> cpu_1f:d_waitrequest
	wire         cpu_1f_data_master_debugaccess;                               // cpu_1f:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1f_data_master_debugaccess
	wire  [18:0] cpu_1f_data_master_address;                                   // cpu_1f:d_address -> mm_interconnect_0:cpu_1f_data_master_address
	wire   [3:0] cpu_1f_data_master_byteenable;                                // cpu_1f:d_byteenable -> mm_interconnect_0:cpu_1f_data_master_byteenable
	wire         cpu_1f_data_master_read;                                      // cpu_1f:d_read -> mm_interconnect_0:cpu_1f_data_master_read
	wire         cpu_1f_data_master_write;                                     // cpu_1f:d_write -> mm_interconnect_0:cpu_1f_data_master_write
	wire  [31:0] cpu_1f_data_master_writedata;                                 // cpu_1f:d_writedata -> mm_interconnect_0:cpu_1f_data_master_writedata
	wire         cpu_1b_p1_mm_bridge_0_m0_waitrequest;                         // mm_interconnect_0:CPU_1b_p1_mm_bridge_0_m0_waitrequest -> CPU_1b_p1:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1b_p1_mm_bridge_0_m0_readdata;                            // mm_interconnect_0:CPU_1b_p1_mm_bridge_0_m0_readdata -> CPU_1b_p1:mm_bridge_0_m0_readdata
	wire         cpu_1b_p1_mm_bridge_0_m0_debugaccess;                         // CPU_1b_p1:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1b_p1_mm_bridge_0_m0_debugaccess
	wire  [16:0] cpu_1b_p1_mm_bridge_0_m0_address;                             // CPU_1b_p1:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1b_p1_mm_bridge_0_m0_address
	wire         cpu_1b_p1_mm_bridge_0_m0_read;                                // CPU_1b_p1:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1b_p1_mm_bridge_0_m0_read
	wire   [3:0] cpu_1b_p1_mm_bridge_0_m0_byteenable;                          // CPU_1b_p1:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1b_p1_mm_bridge_0_m0_byteenable
	wire         cpu_1b_p1_mm_bridge_0_m0_readdatavalid;                       // mm_interconnect_0:CPU_1b_p1_mm_bridge_0_m0_readdatavalid -> CPU_1b_p1:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1b_p1_mm_bridge_0_m0_writedata;                           // CPU_1b_p1:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1b_p1_mm_bridge_0_m0_writedata
	wire         cpu_1b_p1_mm_bridge_0_m0_write;                               // CPU_1b_p1:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1b_p1_mm_bridge_0_m0_write
	wire   [0:0] cpu_1b_p1_mm_bridge_0_m0_burstcount;                          // CPU_1b_p1:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1b_p1_mm_bridge_0_m0_burstcount
	wire         cpu_1e_mm_bridge_0_m0_waitrequest;                            // mm_interconnect_0:CPU_1e_mm_bridge_0_m0_waitrequest -> CPU_1e:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1e_mm_bridge_0_m0_readdata;                               // mm_interconnect_0:CPU_1e_mm_bridge_0_m0_readdata -> CPU_1e:mm_bridge_0_m0_readdata
	wire         cpu_1e_mm_bridge_0_m0_debugaccess;                            // CPU_1e:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_debugaccess
	wire  [16:0] cpu_1e_mm_bridge_0_m0_address;                                // CPU_1e:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_address
	wire         cpu_1e_mm_bridge_0_m0_read;                                   // CPU_1e:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_read
	wire   [3:0] cpu_1e_mm_bridge_0_m0_byteenable;                             // CPU_1e:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_byteenable
	wire         cpu_1e_mm_bridge_0_m0_readdatavalid;                          // mm_interconnect_0:CPU_1e_mm_bridge_0_m0_readdatavalid -> CPU_1e:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1e_mm_bridge_0_m0_writedata;                              // CPU_1e:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_writedata
	wire         cpu_1e_mm_bridge_0_m0_write;                                  // CPU_1e:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_write
	wire   [0:0] cpu_1e_mm_bridge_0_m0_burstcount;                             // CPU_1e:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_burstcount
	wire         cpu_1d_p1_mm_bridge_0_m0_waitrequest;                         // mm_interconnect_0:CPU_1d_p1_mm_bridge_0_m0_waitrequest -> CPU_1d_p1:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1d_p1_mm_bridge_0_m0_readdata;                            // mm_interconnect_0:CPU_1d_p1_mm_bridge_0_m0_readdata -> CPU_1d_p1:mm_bridge_0_m0_readdata
	wire         cpu_1d_p1_mm_bridge_0_m0_debugaccess;                         // CPU_1d_p1:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1d_p1_mm_bridge_0_m0_debugaccess
	wire  [16:0] cpu_1d_p1_mm_bridge_0_m0_address;                             // CPU_1d_p1:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1d_p1_mm_bridge_0_m0_address
	wire         cpu_1d_p1_mm_bridge_0_m0_read;                                // CPU_1d_p1:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1d_p1_mm_bridge_0_m0_read
	wire   [3:0] cpu_1d_p1_mm_bridge_0_m0_byteenable;                          // CPU_1d_p1:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1d_p1_mm_bridge_0_m0_byteenable
	wire         cpu_1d_p1_mm_bridge_0_m0_readdatavalid;                       // mm_interconnect_0:CPU_1d_p1_mm_bridge_0_m0_readdatavalid -> CPU_1d_p1:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1d_p1_mm_bridge_0_m0_writedata;                           // CPU_1d_p1:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1d_p1_mm_bridge_0_m0_writedata
	wire         cpu_1d_p1_mm_bridge_0_m0_write;                               // CPU_1d_p1:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1d_p1_mm_bridge_0_m0_write
	wire   [0:0] cpu_1d_p1_mm_bridge_0_m0_burstcount;                          // CPU_1d_p1:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1d_p1_mm_bridge_0_m0_burstcount
	wire         cpu_1c_p1_mm_bridge_0_m0_waitrequest;                         // mm_interconnect_0:CPU_1c_p1_mm_bridge_0_m0_waitrequest -> CPU_1c_p1:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1c_p1_mm_bridge_0_m0_readdata;                            // mm_interconnect_0:CPU_1c_p1_mm_bridge_0_m0_readdata -> CPU_1c_p1:mm_bridge_0_m0_readdata
	wire         cpu_1c_p1_mm_bridge_0_m0_debugaccess;                         // CPU_1c_p1:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1c_p1_mm_bridge_0_m0_debugaccess
	wire  [16:0] cpu_1c_p1_mm_bridge_0_m0_address;                             // CPU_1c_p1:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1c_p1_mm_bridge_0_m0_address
	wire         cpu_1c_p1_mm_bridge_0_m0_read;                                // CPU_1c_p1:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1c_p1_mm_bridge_0_m0_read
	wire   [3:0] cpu_1c_p1_mm_bridge_0_m0_byteenable;                          // CPU_1c_p1:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1c_p1_mm_bridge_0_m0_byteenable
	wire         cpu_1c_p1_mm_bridge_0_m0_readdatavalid;                       // mm_interconnect_0:CPU_1c_p1_mm_bridge_0_m0_readdatavalid -> CPU_1c_p1:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1c_p1_mm_bridge_0_m0_writedata;                           // CPU_1c_p1:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1c_p1_mm_bridge_0_m0_writedata
	wire         cpu_1c_p1_mm_bridge_0_m0_write;                               // CPU_1c_p1:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1c_p1_mm_bridge_0_m0_write
	wire   [0:0] cpu_1c_p1_mm_bridge_0_m0_burstcount;                          // CPU_1c_p1:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1c_p1_mm_bridge_0_m0_burstcount
	wire         cpu_1b_p2_mm_bridge_0_m0_waitrequest;                         // mm_interconnect_0:CPU_1b_p2_mm_bridge_0_m0_waitrequest -> CPU_1b_p2:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1b_p2_mm_bridge_0_m0_readdata;                            // mm_interconnect_0:CPU_1b_p2_mm_bridge_0_m0_readdata -> CPU_1b_p2:mm_bridge_0_m0_readdata
	wire         cpu_1b_p2_mm_bridge_0_m0_debugaccess;                         // CPU_1b_p2:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1b_p2_mm_bridge_0_m0_debugaccess
	wire  [16:0] cpu_1b_p2_mm_bridge_0_m0_address;                             // CPU_1b_p2:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1b_p2_mm_bridge_0_m0_address
	wire         cpu_1b_p2_mm_bridge_0_m0_read;                                // CPU_1b_p2:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1b_p2_mm_bridge_0_m0_read
	wire   [3:0] cpu_1b_p2_mm_bridge_0_m0_byteenable;                          // CPU_1b_p2:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1b_p2_mm_bridge_0_m0_byteenable
	wire         cpu_1b_p2_mm_bridge_0_m0_readdatavalid;                       // mm_interconnect_0:CPU_1b_p2_mm_bridge_0_m0_readdatavalid -> CPU_1b_p2:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1b_p2_mm_bridge_0_m0_writedata;                           // CPU_1b_p2:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1b_p2_mm_bridge_0_m0_writedata
	wire         cpu_1b_p2_mm_bridge_0_m0_write;                               // CPU_1b_p2:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1b_p2_mm_bridge_0_m0_write
	wire   [0:0] cpu_1b_p2_mm_bridge_0_m0_burstcount;                          // CPU_1b_p2:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1b_p2_mm_bridge_0_m0_burstcount
	wire         cpu_1b_p3_mm_bridge_0_m0_waitrequest;                         // mm_interconnect_0:CPU_1b_p3_mm_bridge_0_m0_waitrequest -> CPU_1b_p3:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1b_p3_mm_bridge_0_m0_readdata;                            // mm_interconnect_0:CPU_1b_p3_mm_bridge_0_m0_readdata -> CPU_1b_p3:mm_bridge_0_m0_readdata
	wire         cpu_1b_p3_mm_bridge_0_m0_debugaccess;                         // CPU_1b_p3:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1b_p3_mm_bridge_0_m0_debugaccess
	wire  [16:0] cpu_1b_p3_mm_bridge_0_m0_address;                             // CPU_1b_p3:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1b_p3_mm_bridge_0_m0_address
	wire         cpu_1b_p3_mm_bridge_0_m0_read;                                // CPU_1b_p3:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1b_p3_mm_bridge_0_m0_read
	wire   [3:0] cpu_1b_p3_mm_bridge_0_m0_byteenable;                          // CPU_1b_p3:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1b_p3_mm_bridge_0_m0_byteenable
	wire         cpu_1b_p3_mm_bridge_0_m0_readdatavalid;                       // mm_interconnect_0:CPU_1b_p3_mm_bridge_0_m0_readdatavalid -> CPU_1b_p3:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1b_p3_mm_bridge_0_m0_writedata;                           // CPU_1b_p3:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1b_p3_mm_bridge_0_m0_writedata
	wire         cpu_1b_p3_mm_bridge_0_m0_write;                               // CPU_1b_p3:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1b_p3_mm_bridge_0_m0_write
	wire   [0:0] cpu_1b_p3_mm_bridge_0_m0_burstcount;                          // CPU_1b_p3:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1b_p3_mm_bridge_0_m0_burstcount
	wire         cpu_1c_p2_mm_bridge_0_m0_waitrequest;                         // mm_interconnect_0:CPU_1c_p2_mm_bridge_0_m0_waitrequest -> CPU_1c_p2:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1c_p2_mm_bridge_0_m0_readdata;                            // mm_interconnect_0:CPU_1c_p2_mm_bridge_0_m0_readdata -> CPU_1c_p2:mm_bridge_0_m0_readdata
	wire         cpu_1c_p2_mm_bridge_0_m0_debugaccess;                         // CPU_1c_p2:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1c_p2_mm_bridge_0_m0_debugaccess
	wire  [16:0] cpu_1c_p2_mm_bridge_0_m0_address;                             // CPU_1c_p2:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1c_p2_mm_bridge_0_m0_address
	wire         cpu_1c_p2_mm_bridge_0_m0_read;                                // CPU_1c_p2:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1c_p2_mm_bridge_0_m0_read
	wire   [3:0] cpu_1c_p2_mm_bridge_0_m0_byteenable;                          // CPU_1c_p2:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1c_p2_mm_bridge_0_m0_byteenable
	wire         cpu_1c_p2_mm_bridge_0_m0_readdatavalid;                       // mm_interconnect_0:CPU_1c_p2_mm_bridge_0_m0_readdatavalid -> CPU_1c_p2:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1c_p2_mm_bridge_0_m0_writedata;                           // CPU_1c_p2:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1c_p2_mm_bridge_0_m0_writedata
	wire         cpu_1c_p2_mm_bridge_0_m0_write;                               // CPU_1c_p2:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1c_p2_mm_bridge_0_m0_write
	wire   [0:0] cpu_1c_p2_mm_bridge_0_m0_burstcount;                          // CPU_1c_p2:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1c_p2_mm_bridge_0_m0_burstcount
	wire         cpu_1c_p3_mm_bridge_0_m0_waitrequest;                         // mm_interconnect_0:CPU_1c_p3_mm_bridge_0_m0_waitrequest -> CPU_1c_p3:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1c_p3_mm_bridge_0_m0_readdata;                            // mm_interconnect_0:CPU_1c_p3_mm_bridge_0_m0_readdata -> CPU_1c_p3:mm_bridge_0_m0_readdata
	wire         cpu_1c_p3_mm_bridge_0_m0_debugaccess;                         // CPU_1c_p3:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1c_p3_mm_bridge_0_m0_debugaccess
	wire  [16:0] cpu_1c_p3_mm_bridge_0_m0_address;                             // CPU_1c_p3:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1c_p3_mm_bridge_0_m0_address
	wire         cpu_1c_p3_mm_bridge_0_m0_read;                                // CPU_1c_p3:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1c_p3_mm_bridge_0_m0_read
	wire   [3:0] cpu_1c_p3_mm_bridge_0_m0_byteenable;                          // CPU_1c_p3:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1c_p3_mm_bridge_0_m0_byteenable
	wire         cpu_1c_p3_mm_bridge_0_m0_readdatavalid;                       // mm_interconnect_0:CPU_1c_p3_mm_bridge_0_m0_readdatavalid -> CPU_1c_p3:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1c_p3_mm_bridge_0_m0_writedata;                           // CPU_1c_p3:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1c_p3_mm_bridge_0_m0_writedata
	wire         cpu_1c_p3_mm_bridge_0_m0_write;                               // CPU_1c_p3:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1c_p3_mm_bridge_0_m0_write
	wire   [0:0] cpu_1c_p3_mm_bridge_0_m0_burstcount;                          // CPU_1c_p3:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1c_p3_mm_bridge_0_m0_burstcount
	wire         cpu_1d_p2_mm_bridge_0_m0_waitrequest;                         // mm_interconnect_0:CPU_1d_p2_mm_bridge_0_m0_waitrequest -> CPU_1d_p2:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1d_p2_mm_bridge_0_m0_readdata;                            // mm_interconnect_0:CPU_1d_p2_mm_bridge_0_m0_readdata -> CPU_1d_p2:mm_bridge_0_m0_readdata
	wire         cpu_1d_p2_mm_bridge_0_m0_debugaccess;                         // CPU_1d_p2:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1d_p2_mm_bridge_0_m0_debugaccess
	wire  [16:0] cpu_1d_p2_mm_bridge_0_m0_address;                             // CPU_1d_p2:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1d_p2_mm_bridge_0_m0_address
	wire         cpu_1d_p2_mm_bridge_0_m0_read;                                // CPU_1d_p2:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1d_p2_mm_bridge_0_m0_read
	wire   [3:0] cpu_1d_p2_mm_bridge_0_m0_byteenable;                          // CPU_1d_p2:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1d_p2_mm_bridge_0_m0_byteenable
	wire         cpu_1d_p2_mm_bridge_0_m0_readdatavalid;                       // mm_interconnect_0:CPU_1d_p2_mm_bridge_0_m0_readdatavalid -> CPU_1d_p2:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1d_p2_mm_bridge_0_m0_writedata;                           // CPU_1d_p2:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1d_p2_mm_bridge_0_m0_writedata
	wire         cpu_1d_p2_mm_bridge_0_m0_write;                               // CPU_1d_p2:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1d_p2_mm_bridge_0_m0_write
	wire   [0:0] cpu_1d_p2_mm_bridge_0_m0_burstcount;                          // CPU_1d_p2:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1d_p2_mm_bridge_0_m0_burstcount
	wire         cpu_1d_p3_mm_bridge_0_m0_waitrequest;                         // mm_interconnect_0:CPU_1d_p3_mm_bridge_0_m0_waitrequest -> CPU_1d_p3:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1d_p3_mm_bridge_0_m0_readdata;                            // mm_interconnect_0:CPU_1d_p3_mm_bridge_0_m0_readdata -> CPU_1d_p3:mm_bridge_0_m0_readdata
	wire         cpu_1d_p3_mm_bridge_0_m0_debugaccess;                         // CPU_1d_p3:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1d_p3_mm_bridge_0_m0_debugaccess
	wire  [16:0] cpu_1d_p3_mm_bridge_0_m0_address;                             // CPU_1d_p3:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1d_p3_mm_bridge_0_m0_address
	wire         cpu_1d_p3_mm_bridge_0_m0_read;                                // CPU_1d_p3:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1d_p3_mm_bridge_0_m0_read
	wire   [3:0] cpu_1d_p3_mm_bridge_0_m0_byteenable;                          // CPU_1d_p3:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1d_p3_mm_bridge_0_m0_byteenable
	wire         cpu_1d_p3_mm_bridge_0_m0_readdatavalid;                       // mm_interconnect_0:CPU_1d_p3_mm_bridge_0_m0_readdatavalid -> CPU_1d_p3:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1d_p3_mm_bridge_0_m0_writedata;                           // CPU_1d_p3:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1d_p3_mm_bridge_0_m0_writedata
	wire         cpu_1d_p3_mm_bridge_0_m0_write;                               // CPU_1d_p3:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1d_p3_mm_bridge_0_m0_write
	wire   [0:0] cpu_1d_p3_mm_bridge_0_m0_burstcount;                          // CPU_1d_p3:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1d_p3_mm_bridge_0_m0_burstcount
	wire  [31:0] cpu_1f_instruction_master_readdata;                           // mm_interconnect_0:cpu_1f_instruction_master_readdata -> cpu_1f:i_readdata
	wire         cpu_1f_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_1f_instruction_master_waitrequest -> cpu_1f:i_waitrequest
	wire  [18:0] cpu_1f_instruction_master_address;                            // cpu_1f:i_address -> mm_interconnect_0:cpu_1f_instruction_master_address
	wire         cpu_1f_instruction_master_read;                               // cpu_1f:i_read -> mm_interconnect_0:cpu_1f_instruction_master_read
	wire  [31:0] cpu_1a_instruction_master_readdata;                           // mm_interconnect_0:cpu_1a_instruction_master_readdata -> cpu_1a:i_readdata
	wire         cpu_1a_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_1a_instruction_master_waitrequest -> cpu_1a:i_waitrequest
	wire  [27:0] cpu_1a_instruction_master_address;                            // cpu_1a:i_address -> mm_interconnect_0:cpu_1a_instruction_master_address
	wire         cpu_1a_instruction_master_read;                               // cpu_1a:i_read -> mm_interconnect_0:cpu_1a_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1a_avalon_jtag_slave_chipselect -> jtag_uart_1a:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_readdata;    // jtag_uart_1a:av_readdata -> mm_interconnect_0:jtag_uart_1a_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_waitrequest; // jtag_uart_1a:av_waitrequest -> mm_interconnect_0:jtag_uart_1a_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1a_avalon_jtag_slave_address -> jtag_uart_1a:av_address
	wire         mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1a_avalon_jtag_slave_read -> jtag_uart_1a:av_read_n
	wire         mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1a_avalon_jtag_slave_write -> jtag_uart_1a:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1a_avalon_jtag_slave_writedata -> jtag_uart_1a:av_writedata
	wire  [31:0] mm_interconnect_0_sys_id_1a_control_slave_readdata;           // sys_id_1a:readdata -> mm_interconnect_0:sys_id_1a_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sys_id_1a_control_slave_address;            // mm_interconnect_0:sys_id_1a_control_slave_address -> sys_id_1a:address
	wire  [31:0] mm_interconnect_0_cpu_1a_debug_mem_slave_readdata;            // cpu_1a:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1a_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_1a_debug_mem_slave_waitrequest;         // cpu_1a:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1a_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_1a_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_1a_debug_mem_slave_debugaccess -> cpu_1a:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_1a_debug_mem_slave_address;             // mm_interconnect_0:cpu_1a_debug_mem_slave_address -> cpu_1a:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_1a_debug_mem_slave_read;                // mm_interconnect_0:cpu_1a_debug_mem_slave_read -> cpu_1a:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_1a_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_1a_debug_mem_slave_byteenable -> cpu_1a:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_1a_debug_mem_slave_write;               // mm_interconnect_0:cpu_1a_debug_mem_slave_write -> cpu_1a:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_1a_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_1a_debug_mem_slave_writedata -> cpu_1a:debug_mem_slave_writedata
	wire         mm_interconnect_0_fifo_qa_p1_in_waitrequest;                  // fifo_qa_p1:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qa_p1_in_waitrequest
	wire         mm_interconnect_0_fifo_qa_p1_in_write;                        // mm_interconnect_0:fifo_qa_p1_in_write -> fifo_qa_p1:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qa_p1_in_writedata;                    // mm_interconnect_0:fifo_qa_p1_in_writedata -> fifo_qa_p1:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_qa_p2_in_waitrequest;                  // fifo_qa_p2:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qa_p2_in_waitrequest
	wire         mm_interconnect_0_fifo_qa_p2_in_write;                        // mm_interconnect_0:fifo_qa_p2_in_write -> fifo_qa_p2:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qa_p2_in_writedata;                    // mm_interconnect_0:fifo_qa_p2_in_writedata -> fifo_qa_p2:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_qa_p3_in_waitrequest;                  // fifo_qa_p3:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qa_p3_in_waitrequest
	wire         mm_interconnect_0_fifo_qa_p3_in_write;                        // mm_interconnect_0:fifo_qa_p3_in_write -> fifo_qa_p3:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qa_p3_in_writedata;                    // mm_interconnect_0:fifo_qa_p3_in_writedata -> fifo_qa_p3:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qa_p1_in_csr_readdata;                 // fifo_qa_p1:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qa_p1_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qa_p1_in_csr_address;                  // mm_interconnect_0:fifo_qa_p1_in_csr_address -> fifo_qa_p1:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qa_p1_in_csr_read;                     // mm_interconnect_0:fifo_qa_p1_in_csr_read -> fifo_qa_p1:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qa_p1_in_csr_write;                    // mm_interconnect_0:fifo_qa_p1_in_csr_write -> fifo_qa_p1:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qa_p1_in_csr_writedata;                // mm_interconnect_0:fifo_qa_p1_in_csr_writedata -> fifo_qa_p1:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qa_p2_in_csr_readdata;                 // fifo_qa_p2:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qa_p2_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qa_p2_in_csr_address;                  // mm_interconnect_0:fifo_qa_p2_in_csr_address -> fifo_qa_p2:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qa_p2_in_csr_read;                     // mm_interconnect_0:fifo_qa_p2_in_csr_read -> fifo_qa_p2:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qa_p2_in_csr_write;                    // mm_interconnect_0:fifo_qa_p2_in_csr_write -> fifo_qa_p2:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qa_p2_in_csr_writedata;                // mm_interconnect_0:fifo_qa_p2_in_csr_writedata -> fifo_qa_p2:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qa_p3_in_csr_readdata;                 // fifo_qa_p3:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qa_p3_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qa_p3_in_csr_address;                  // mm_interconnect_0:fifo_qa_p3_in_csr_address -> fifo_qa_p3:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qa_p3_in_csr_read;                     // mm_interconnect_0:fifo_qa_p3_in_csr_read -> fifo_qa_p3:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qa_p3_in_csr_write;                    // mm_interconnect_0:fifo_qa_p3_in_csr_write -> fifo_qa_p3:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qa_p3_in_csr_writedata;                // mm_interconnect_0:fifo_qa_p3_in_csr_writedata -> fifo_qa_p3:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                     // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                      // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                         // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                        // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                    // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;             // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;               // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;            // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;                // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;                   // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;             // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;          // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;                  // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;              // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         mm_interconnect_0_timer_1a_s1_chipselect;                     // mm_interconnect_0:timer_1a_s1_chipselect -> timer_1a:chipselect
	wire  [15:0] mm_interconnect_0_timer_1a_s1_readdata;                       // timer_1a:readdata -> mm_interconnect_0:timer_1a_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1a_s1_address;                        // mm_interconnect_0:timer_1a_s1_address -> timer_1a:address
	wire         mm_interconnect_0_timer_1a_s1_write;                          // mm_interconnect_0:timer_1a_s1_write -> timer_1a:write_n
	wire  [15:0] mm_interconnect_0_timer_1a_s1_writedata;                      // mm_interconnect_0:timer_1a_s1_writedata -> timer_1a:writedata
	wire         mm_interconnect_0_mem_info_s1_chipselect;                     // mm_interconnect_0:mem_info_s1_chipselect -> mem_info:chipselect
	wire  [31:0] mm_interconnect_0_mem_info_s1_readdata;                       // mem_info:readdata -> mm_interconnect_0:mem_info_s1_readdata
	wire   [7:0] mm_interconnect_0_mem_info_s1_address;                        // mm_interconnect_0:mem_info_s1_address -> mem_info:address
	wire   [3:0] mm_interconnect_0_mem_info_s1_byteenable;                     // mm_interconnect_0:mem_info_s1_byteenable -> mem_info:byteenable
	wire         mm_interconnect_0_mem_info_s1_write;                          // mm_interconnect_0:mem_info_s1_write -> mem_info:write
	wire  [31:0] mm_interconnect_0_mem_info_s1_writedata;                      // mm_interconnect_0:mem_info_s1_writedata -> mem_info:writedata
	wire         mm_interconnect_0_mem_info_s1_clken;                          // mm_interconnect_0:mem_info_s1_clken -> mem_info:clken
	wire         mm_interconnect_0_fifo_qd_p3_in_waitrequest;                  // fifo_qd_p3:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qd_p3_in_waitrequest
	wire         mm_interconnect_0_fifo_qd_p3_in_write;                        // mm_interconnect_0:fifo_qd_p3_in_write -> fifo_qd_p3:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qd_p3_in_writedata;                    // mm_interconnect_0:fifo_qd_p3_in_writedata -> fifo_qd_p3:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qc_p3_in_csr_readdata;                 // fifo_qc_p3:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qc_p3_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qc_p3_in_csr_address;                  // mm_interconnect_0:fifo_qc_p3_in_csr_address -> fifo_qc_p3:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qc_p3_in_csr_read;                     // mm_interconnect_0:fifo_qc_p3_in_csr_read -> fifo_qc_p3:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qc_p3_in_csr_write;                    // mm_interconnect_0:fifo_qc_p3_in_csr_write -> fifo_qc_p3:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qc_p3_in_csr_writedata;                // mm_interconnect_0:fifo_qc_p3_in_csr_writedata -> fifo_qc_p3:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qd_p3_in_csr_readdata;                 // fifo_qd_p3:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qd_p3_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qd_p3_in_csr_address;                  // mm_interconnect_0:fifo_qd_p3_in_csr_address -> fifo_qd_p3:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qd_p3_in_csr_read;                     // mm_interconnect_0:fifo_qd_p3_in_csr_read -> fifo_qd_p3:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qd_p3_in_csr_write;                    // mm_interconnect_0:fifo_qd_p3_in_csr_write -> fifo_qd_p3:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qd_p3_in_csr_writedata;                // mm_interconnect_0:fifo_qd_p3_in_csr_writedata -> fifo_qd_p3:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qc_p3_out_readdata;                    // fifo_qc_p3:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qc_p3_out_readdata
	wire         mm_interconnect_0_fifo_qc_p3_out_waitrequest;                 // fifo_qc_p3:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qc_p3_out_waitrequest
	wire         mm_interconnect_0_fifo_qc_p3_out_read;                        // mm_interconnect_0:fifo_qc_p3_out_read -> fifo_qc_p3:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_qe_in_waitrequest;                     // fifo_qe:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qe_in_waitrequest
	wire         mm_interconnect_0_fifo_qe_in_write;                           // mm_interconnect_0:fifo_qe_in_write -> fifo_qe:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qe_in_writedata;                       // mm_interconnect_0:fifo_qe_in_writedata -> fifo_qe:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qd_p1_in_csr_readdata;                 // fifo_qd_p1:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qd_p1_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qd_p1_in_csr_address;                  // mm_interconnect_0:fifo_qd_p1_in_csr_address -> fifo_qd_p1:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qd_p1_in_csr_read;                     // mm_interconnect_0:fifo_qd_p1_in_csr_read -> fifo_qd_p1:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qd_p1_in_csr_write;                    // mm_interconnect_0:fifo_qd_p1_in_csr_write -> fifo_qd_p1:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qd_p1_in_csr_writedata;                // mm_interconnect_0:fifo_qd_p1_in_csr_writedata -> fifo_qd_p1:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qe_in_csr_readdata;                    // fifo_qe:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qe_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qe_in_csr_address;                     // mm_interconnect_0:fifo_qe_in_csr_address -> fifo_qe:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qe_in_csr_read;                        // mm_interconnect_0:fifo_qe_in_csr_read -> fifo_qe:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qe_in_csr_write;                       // mm_interconnect_0:fifo_qe_in_csr_write -> fifo_qe:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qe_in_csr_writedata;                   // mm_interconnect_0:fifo_qe_in_csr_writedata -> fifo_qe:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qd_p2_in_csr_readdata;                 // fifo_qd_p2:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qd_p2_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qd_p2_in_csr_address;                  // mm_interconnect_0:fifo_qd_p2_in_csr_address -> fifo_qd_p2:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qd_p2_in_csr_read;                     // mm_interconnect_0:fifo_qd_p2_in_csr_read -> fifo_qd_p2:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qd_p2_in_csr_write;                    // mm_interconnect_0:fifo_qd_p2_in_csr_write -> fifo_qd_p2:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qd_p2_in_csr_writedata;                // mm_interconnect_0:fifo_qd_p2_in_csr_writedata -> fifo_qd_p2:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qd_p1_out_readdata;                    // fifo_qd_p1:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qd_p1_out_readdata
	wire         mm_interconnect_0_fifo_qd_p1_out_waitrequest;                 // fifo_qd_p1:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qd_p1_out_waitrequest
	wire         mm_interconnect_0_fifo_qd_p1_out_read;                        // mm_interconnect_0:fifo_qd_p1_out_read -> fifo_qd_p1:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_qd_p2_out_readdata;                    // fifo_qd_p2:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qd_p2_out_readdata
	wire         mm_interconnect_0_fifo_qd_p2_out_waitrequest;                 // fifo_qd_p2:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qd_p2_out_waitrequest
	wire         mm_interconnect_0_fifo_qd_p2_out_read;                        // mm_interconnect_0:fifo_qd_p2_out_read -> fifo_qd_p2:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_qd_p3_out_readdata;                    // fifo_qd_p3:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qd_p3_out_readdata
	wire         mm_interconnect_0_fifo_qd_p3_out_waitrequest;                 // fifo_qd_p3:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qd_p3_out_waitrequest
	wire         mm_interconnect_0_fifo_qd_p3_out_read;                        // mm_interconnect_0:fifo_qd_p3_out_read -> fifo_qd_p3:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_qd_p2_in_waitrequest;                  // fifo_qd_p2:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qd_p2_in_waitrequest
	wire         mm_interconnect_0_fifo_qd_p2_in_write;                        // mm_interconnect_0:fifo_qd_p2_in_write -> fifo_qd_p2:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qd_p2_in_writedata;                    // mm_interconnect_0:fifo_qd_p2_in_writedata -> fifo_qd_p2:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qc_p2_in_csr_readdata;                 // fifo_qc_p2:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qc_p2_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qc_p2_in_csr_address;                  // mm_interconnect_0:fifo_qc_p2_in_csr_address -> fifo_qc_p2:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qc_p2_in_csr_read;                     // mm_interconnect_0:fifo_qc_p2_in_csr_read -> fifo_qc_p2:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qc_p2_in_csr_write;                    // mm_interconnect_0:fifo_qc_p2_in_csr_write -> fifo_qc_p2:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qc_p2_in_csr_writedata;                // mm_interconnect_0:fifo_qc_p2_in_csr_writedata -> fifo_qc_p2:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qc_p2_out_readdata;                    // fifo_qc_p2:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qc_p2_out_readdata
	wire         mm_interconnect_0_fifo_qc_p2_out_waitrequest;                 // fifo_qc_p2:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qc_p2_out_waitrequest
	wire         mm_interconnect_0_fifo_qc_p2_out_read;                        // mm_interconnect_0:fifo_qc_p2_out_read -> fifo_qc_p2:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_qc_p2_in_waitrequest;                  // fifo_qc_p2:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qc_p2_in_waitrequest
	wire         mm_interconnect_0_fifo_qc_p2_in_write;                        // mm_interconnect_0:fifo_qc_p2_in_write -> fifo_qc_p2:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qc_p2_in_writedata;                    // mm_interconnect_0:fifo_qc_p2_in_writedata -> fifo_qc_p2:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qb_p2_in_csr_readdata;                 // fifo_qb_p2:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qb_p2_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qb_p2_in_csr_address;                  // mm_interconnect_0:fifo_qb_p2_in_csr_address -> fifo_qb_p2:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qb_p2_in_csr_read;                     // mm_interconnect_0:fifo_qb_p2_in_csr_read -> fifo_qb_p2:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qb_p2_in_csr_write;                    // mm_interconnect_0:fifo_qb_p2_in_csr_write -> fifo_qb_p2:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qb_p2_in_csr_writedata;                // mm_interconnect_0:fifo_qb_p2_in_csr_writedata -> fifo_qb_p2:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qb_p2_out_readdata;                    // fifo_qb_p2:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qb_p2_out_readdata
	wire         mm_interconnect_0_fifo_qb_p2_out_waitrequest;                 // fifo_qb_p2:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qb_p2_out_waitrequest
	wire         mm_interconnect_0_fifo_qb_p2_out_read;                        // mm_interconnect_0:fifo_qb_p2_out_read -> fifo_qb_p2:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_qb_p2_in_waitrequest;                  // fifo_qb_p2:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qb_p2_in_waitrequest
	wire         mm_interconnect_0_fifo_qb_p2_in_write;                        // mm_interconnect_0:fifo_qb_p2_in_write -> fifo_qb_p2:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qb_p2_in_writedata;                    // mm_interconnect_0:fifo_qb_p2_in_writedata -> fifo_qb_p2:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qa_p2_out_readdata;                    // fifo_qa_p2:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qa_p2_out_readdata
	wire         mm_interconnect_0_fifo_qa_p2_out_waitrequest;                 // fifo_qa_p2:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qa_p2_out_waitrequest
	wire         mm_interconnect_0_fifo_qa_p2_out_read;                        // mm_interconnect_0:fifo_qa_p2_out_read -> fifo_qa_p2:avalonmm_read_slave_read
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_chipselect -> jtag_uart_1f:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_readdata;    // jtag_uart_1f:av_readdata -> mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_waitrequest; // jtag_uart_1f:av_waitrequest -> mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_address -> jtag_uart_1f:av_address
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_read -> jtag_uart_1f:av_read_n
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_write -> jtag_uart_1f:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_writedata -> jtag_uart_1f:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_1f_control_slave_readdata;            // sysid_1f:readdata -> mm_interconnect_0:sysid_1f_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_1f_control_slave_address;             // mm_interconnect_0:sysid_1f_control_slave_address -> sysid_1f:address
	wire  [31:0] mm_interconnect_0_cpu_1f_debug_mem_slave_readdata;            // cpu_1f:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1f_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_1f_debug_mem_slave_waitrequest;         // cpu_1f:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1f_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_1f_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_1f_debug_mem_slave_debugaccess -> cpu_1f:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_1f_debug_mem_slave_address;             // mm_interconnect_0:cpu_1f_debug_mem_slave_address -> cpu_1f:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_1f_debug_mem_slave_read;                // mm_interconnect_0:cpu_1f_debug_mem_slave_read -> cpu_1f:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_1f_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_1f_debug_mem_slave_byteenable -> cpu_1f:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_1f_debug_mem_slave_write;               // mm_interconnect_0:cpu_1f_debug_mem_slave_write -> cpu_1f:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_1f_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_1f_debug_mem_slave_writedata -> cpu_1f:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qe_out_readdata;                       // fifo_qe:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qe_out_readdata
	wire         mm_interconnect_0_fifo_qe_out_waitrequest;                    // fifo_qe:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qe_out_waitrequest
	wire         mm_interconnect_0_fifo_qe_out_read;                           // mm_interconnect_0:fifo_qe_out_read -> fifo_qe:avalonmm_read_slave_read
	wire         mm_interconnect_0_timer_1f_s1_chipselect;                     // mm_interconnect_0:timer_1f_s1_chipselect -> timer_1f:chipselect
	wire  [15:0] mm_interconnect_0_timer_1f_s1_readdata;                       // timer_1f:readdata -> mm_interconnect_0:timer_1f_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1f_s1_address;                        // mm_interconnect_0:timer_1f_s1_address -> timer_1f:address
	wire         mm_interconnect_0_timer_1f_s1_write;                          // mm_interconnect_0:timer_1f_s1_write -> timer_1f:write_n
	wire  [15:0] mm_interconnect_0_timer_1f_s1_writedata;                      // mm_interconnect_0:timer_1f_s1_writedata -> timer_1f:writedata
	wire         mm_interconnect_0_oc_ram_1f_s1_chipselect;                    // mm_interconnect_0:oc_ram_1f_s1_chipselect -> oc_ram_1f:chipselect
	wire  [31:0] mm_interconnect_0_oc_ram_1f_s1_readdata;                      // oc_ram_1f:readdata -> mm_interconnect_0:oc_ram_1f_s1_readdata
	wire  [14:0] mm_interconnect_0_oc_ram_1f_s1_address;                       // mm_interconnect_0:oc_ram_1f_s1_address -> oc_ram_1f:address
	wire   [3:0] mm_interconnect_0_oc_ram_1f_s1_byteenable;                    // mm_interconnect_0:oc_ram_1f_s1_byteenable -> oc_ram_1f:byteenable
	wire         mm_interconnect_0_oc_ram_1f_s1_write;                         // mm_interconnect_0:oc_ram_1f_s1_write -> oc_ram_1f:write
	wire  [31:0] mm_interconnect_0_oc_ram_1f_s1_writedata;                     // mm_interconnect_0:oc_ram_1f_s1_writedata -> oc_ram_1f:writedata
	wire         mm_interconnect_0_oc_ram_1f_s1_clken;                         // mm_interconnect_0:oc_ram_1f_s1_clken -> oc_ram_1f:clken
	wire         mm_interconnect_0_fifo_qd_p1_in_waitrequest;                  // fifo_qd_p1:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qd_p1_in_waitrequest
	wire         mm_interconnect_0_fifo_qd_p1_in_write;                        // mm_interconnect_0:fifo_qd_p1_in_write -> fifo_qd_p1:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qd_p1_in_writedata;                    // mm_interconnect_0:fifo_qd_p1_in_writedata -> fifo_qd_p1:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qc_p1_in_csr_readdata;                 // fifo_qc_p1:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qc_p1_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qc_p1_in_csr_address;                  // mm_interconnect_0:fifo_qc_p1_in_csr_address -> fifo_qc_p1:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qc_p1_in_csr_read;                     // mm_interconnect_0:fifo_qc_p1_in_csr_read -> fifo_qc_p1:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qc_p1_in_csr_write;                    // mm_interconnect_0:fifo_qc_p1_in_csr_write -> fifo_qc_p1:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qc_p1_in_csr_writedata;                // mm_interconnect_0:fifo_qc_p1_in_csr_writedata -> fifo_qc_p1:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qc_p1_out_readdata;                    // fifo_qc_p1:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qc_p1_out_readdata
	wire         mm_interconnect_0_fifo_qc_p1_out_waitrequest;                 // fifo_qc_p1:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qc_p1_out_waitrequest
	wire         mm_interconnect_0_fifo_qc_p1_out_read;                        // mm_interconnect_0:fifo_qc_p1_out_read -> fifo_qc_p1:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_qc_p1_in_waitrequest;                  // fifo_qc_p1:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qc_p1_in_waitrequest
	wire         mm_interconnect_0_fifo_qc_p1_in_write;                        // mm_interconnect_0:fifo_qc_p1_in_write -> fifo_qc_p1:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qc_p1_in_writedata;                    // mm_interconnect_0:fifo_qc_p1_in_writedata -> fifo_qc_p1:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qb_p1_in_csr_readdata;                 // fifo_qb_p1:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qb_p1_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qb_p1_in_csr_address;                  // mm_interconnect_0:fifo_qb_p1_in_csr_address -> fifo_qb_p1:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qb_p1_in_csr_read;                     // mm_interconnect_0:fifo_qb_p1_in_csr_read -> fifo_qb_p1:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qb_p1_in_csr_write;                    // mm_interconnect_0:fifo_qb_p1_in_csr_write -> fifo_qb_p1:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qb_p1_in_csr_writedata;                // mm_interconnect_0:fifo_qb_p1_in_csr_writedata -> fifo_qb_p1:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qb_p1_out_readdata;                    // fifo_qb_p1:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qb_p1_out_readdata
	wire         mm_interconnect_0_fifo_qb_p1_out_waitrequest;                 // fifo_qb_p1:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qb_p1_out_waitrequest
	wire         mm_interconnect_0_fifo_qb_p1_out_read;                        // mm_interconnect_0:fifo_qb_p1_out_read -> fifo_qb_p1:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_qb_p1_in_waitrequest;                  // fifo_qb_p1:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qb_p1_in_waitrequest
	wire         mm_interconnect_0_fifo_qb_p1_in_write;                        // mm_interconnect_0:fifo_qb_p1_in_write -> fifo_qb_p1:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qb_p1_in_writedata;                    // mm_interconnect_0:fifo_qb_p1_in_writedata -> fifo_qb_p1:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qa_p1_out_readdata;                    // fifo_qa_p1:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qa_p1_out_readdata
	wire         mm_interconnect_0_fifo_qa_p1_out_waitrequest;                 // fifo_qa_p1:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qa_p1_out_waitrequest
	wire         mm_interconnect_0_fifo_qa_p1_out_read;                        // mm_interconnect_0:fifo_qa_p1_out_read -> fifo_qa_p1:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_qc_p3_in_waitrequest;                  // fifo_qc_p3:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qc_p3_in_waitrequest
	wire         mm_interconnect_0_fifo_qc_p3_in_write;                        // mm_interconnect_0:fifo_qc_p3_in_write -> fifo_qc_p3:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qc_p3_in_writedata;                    // mm_interconnect_0:fifo_qc_p3_in_writedata -> fifo_qc_p3:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qb_p3_in_csr_readdata;                 // fifo_qb_p3:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_qb_p3_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_qb_p3_in_csr_address;                  // mm_interconnect_0:fifo_qb_p3_in_csr_address -> fifo_qb_p3:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_qb_p3_in_csr_read;                     // mm_interconnect_0:fifo_qb_p3_in_csr_read -> fifo_qb_p3:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_qb_p3_in_csr_write;                    // mm_interconnect_0:fifo_qb_p3_in_csr_write -> fifo_qb_p3:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qb_p3_in_csr_writedata;                // mm_interconnect_0:fifo_qb_p3_in_csr_writedata -> fifo_qb_p3:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qb_p3_out_readdata;                    // fifo_qb_p3:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qb_p3_out_readdata
	wire         mm_interconnect_0_fifo_qb_p3_out_waitrequest;                 // fifo_qb_p3:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qb_p3_out_waitrequest
	wire         mm_interconnect_0_fifo_qb_p3_out_read;                        // mm_interconnect_0:fifo_qb_p3_out_read -> fifo_qb_p3:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_qb_p3_in_waitrequest;                  // fifo_qb_p3:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_qb_p3_in_waitrequest
	wire         mm_interconnect_0_fifo_qb_p3_in_write;                        // mm_interconnect_0:fifo_qb_p3_in_write -> fifo_qb_p3:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_qb_p3_in_writedata;                    // mm_interconnect_0:fifo_qb_p3_in_writedata -> fifo_qb_p3:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_qa_p3_out_readdata;                    // fifo_qa_p3:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_qa_p3_out_readdata
	wire         mm_interconnect_0_fifo_qa_p3_out_waitrequest;                 // fifo_qa_p3:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_qa_p3_out_waitrequest
	wire         mm_interconnect_0_fifo_qa_p3_out_read;                        // mm_interconnect_0:fifo_qa_p3_out_read -> fifo_qa_p3:avalonmm_read_slave_read
	wire         irq_mapper_receiver0_irq;                                     // timer_1a:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart_1a:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_1a_irq_irq;                                               // irq_mapper:sender_irq -> cpu_1a:irq
	wire         irq_mapper_001_receiver0_irq;                                 // timer_1f:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                 // jtag_uart_1f:av_irq -> irq_mapper_001:receiver1_irq
	wire  [31:0] cpu_1f_irq_irq;                                               // irq_mapper_001:sender_irq -> cpu_1f:irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [CPU_1b_p1:reset_bridge_0_in_reset_reset, CPU_1b_p2:reset_bridge_0_in_reset_reset, CPU_1b_p3:reset_bridge_0_in_reset_reset, CPU_1c_p1:reset_bridge_0_in_reset_reset, CPU_1c_p2:reset_bridge_0_in_reset_reset, CPU_1c_p3:reset_bridge_0_in_reset_reset, CPU_1d_p1:reset_bridge_0_in_reset_reset, CPU_1d_p2:reset_bridge_0_in_reset_reset, CPU_1d_p3:reset_bridge_0_in_reset_reset, CPU_1e:reset_bridge_0_in_reset_reset, cpu_1a:reset_n, cpu_1f:reset_n, fifo_qa_p1:reset_n, fifo_qa_p2:reset_n, fifo_qa_p3:reset_n, fifo_qb_p1:reset_n, fifo_qb_p2:reset_n, fifo_qb_p3:reset_n, fifo_qc_p1:reset_n, fifo_qc_p2:reset_n, fifo_qc_p3:reset_n, fifo_qd_p1:reset_n, fifo_qd_p2:reset_n, fifo_qd_p3:reset_n, fifo_qe:reset_n, irq_mapper:reset, irq_mapper_001:reset, jtag_uart_1a:rst_n, jtag_uart_1f:rst_n, mem_info:reset, mm_interconnect_0:cpu_1a_reset_reset_bridge_in_reset_reset, oc_ram_1f:reset, rst_translator:in_reset, sdram_controller:reset_n, sys_id_1a:reset_n, sysid_1f:reset_n, timer_1a:reset_n, timer_1f:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [cpu_1a:reset_req, cpu_1f:reset_req, mem_info:reset_req, oc_ram_1f:reset_req, rst_translator:reset_req_in]
	wire         cpu_1a_debug_reset_request_reset;                             // cpu_1a:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         cpu_1f_debug_reset_request_reset;                             // cpu_1f:debug_reset_request -> [rst_controller:reset_in2, rst_controller_001:reset_in2]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	FTOP_MSOC_CPU_1b_p1 cpu_1b_p1 (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                             //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1b_p1_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1b_p1_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1b_p1_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1b_p1_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1b_p1_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1b_p1_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1b_p1_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1b_p1_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1b_p1_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1b_p1_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)          // reset_bridge_0_in_reset.reset
	);

	FTOP_MSOC_CPU_1b_p2 cpu_1b_p2 (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                             //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1b_p2_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1b_p2_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1b_p2_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1b_p2_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1b_p2_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1b_p2_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1b_p2_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1b_p2_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1b_p2_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1b_p2_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)          // reset_bridge_0_in_reset.reset
	);

	FTOP_MSOC_CPU_1b_p3 cpu_1b_p3 (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                             //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1b_p3_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1b_p3_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1b_p3_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1b_p3_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1b_p3_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1b_p3_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1b_p3_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1b_p3_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1b_p3_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1b_p3_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)          // reset_bridge_0_in_reset.reset
	);

	FTOP_MSOC_CPU_1c_p1 cpu_1c_p1 (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                             //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1c_p1_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1c_p1_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1c_p1_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1c_p1_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1c_p1_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1c_p1_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1c_p1_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1c_p1_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1c_p1_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1c_p1_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)          // reset_bridge_0_in_reset.reset
	);

	FTOP_MSOC_CPU_1c_p2 cpu_1c_p2 (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                             //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1c_p2_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1c_p2_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1c_p2_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1c_p2_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1c_p2_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1c_p2_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1c_p2_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1c_p2_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1c_p2_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1c_p2_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)          // reset_bridge_0_in_reset.reset
	);

	FTOP_MSOC_CPU_1c_p3 cpu_1c_p3 (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                             //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1c_p3_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1c_p3_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1c_p3_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1c_p3_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1c_p3_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1c_p3_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1c_p3_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1c_p3_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1c_p3_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1c_p3_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)          // reset_bridge_0_in_reset.reset
	);

	FTOP_MSOC_CPU_1d_p1 cpu_1d_p1 (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                             //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1d_p1_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1d_p1_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1d_p1_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1d_p1_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1d_p1_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1d_p1_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1d_p1_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1d_p1_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1d_p1_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1d_p1_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)          // reset_bridge_0_in_reset.reset
	);

	FTOP_MSOC_CPU_1d_p2 cpu_1d_p2 (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                             //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1d_p2_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1d_p2_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1d_p2_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1d_p2_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1d_p2_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1d_p2_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1d_p2_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1d_p2_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1d_p2_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1d_p2_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)          // reset_bridge_0_in_reset.reset
	);

	FTOP_MSOC_CPU_1d_p3 cpu_1d_p3 (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                             //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1d_p3_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1d_p3_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1d_p3_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1d_p3_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1d_p3_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1d_p3_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1d_p3_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1d_p3_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1d_p3_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1d_p3_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)          // reset_bridge_0_in_reset.reset
	);

	FTOP_MSOC_CPU_1e cpu_1e (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                          //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1e_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1e_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1e_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1e_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1e_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1e_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1e_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1e_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1e_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1e_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)       // reset_bridge_0_in_reset.reset
	);

	FTOP_MSOC_cpu_1a cpu_1a (
		.clk                                 (pll_c0_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (cpu_1a_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_1a_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_1a_data_master_read),                              //                          .read
		.d_readdata                          (cpu_1a_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_1a_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_1a_data_master_write),                             //                          .write
		.d_writedata                         (cpu_1a_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_1a_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_1a_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_1a_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_1a_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_1a_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_1a_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_1a_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_1a_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_1a_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_1a_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_1a_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_1a_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_1a_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_1a_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_1a_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	FTOP_MSOC_cpu_1f cpu_1f (
		.clk                                 (pll_c0_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (cpu_1f_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_1f_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_1f_data_master_read),                              //                          .read
		.d_readdata                          (cpu_1f_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_1f_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_1f_data_master_write),                             //                          .write
		.d_writedata                         (cpu_1f_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_1f_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_1f_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_1f_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_1f_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_1f_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_1f_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_1f_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_1f_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_1f_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_1f_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_1f_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_1f_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_1f_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_1f_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_1f_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	FTOP_MSOC_fifo_qa_p1 fifo_qa_p1 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qa_p1_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qa_p1_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qa_p1_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qa_p1_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qa_p1_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qa_p1_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qa_p1_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qa_p1_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qa_p1_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qa_p1_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qa_p1_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qa_p1 fifo_qa_p2 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qa_p2_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qa_p2_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qa_p2_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qa_p2_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qa_p2_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qa_p2_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qa_p2_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qa_p2_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qa_p2_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qa_p2_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qa_p2_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qa_p1 fifo_qa_p3 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qa_p3_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qa_p3_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qa_p3_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qa_p3_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qa_p3_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qa_p3_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qa_p3_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qa_p3_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qa_p3_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qa_p3_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qa_p3_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qb_p1 fifo_qb_p1 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qb_p1_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qb_p1_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qb_p1_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qb_p1_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qb_p1_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qb_p1_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qb_p1_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qb_p1_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qb_p1_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qb_p1_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qb_p1_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qb_p1 fifo_qb_p2 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qb_p2_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qb_p2_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qb_p2_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qb_p2_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qb_p2_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qb_p2_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qb_p2_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qb_p2_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qb_p2_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qb_p2_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qb_p2_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qb_p1 fifo_qb_p3 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qb_p3_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qb_p3_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qb_p3_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qb_p3_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qb_p3_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qb_p3_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qb_p3_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qb_p3_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qb_p3_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qb_p3_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qb_p3_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qb_p1 fifo_qc_p1 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qc_p1_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qc_p1_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qc_p1_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qc_p1_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qc_p1_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qc_p1_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qc_p1_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qc_p1_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qc_p1_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qc_p1_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qc_p1_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qb_p1 fifo_qc_p2 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qc_p2_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qc_p2_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qc_p2_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qc_p2_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qc_p2_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qc_p2_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qc_p2_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qc_p2_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qc_p2_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qc_p2_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qc_p2_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qb_p1 fifo_qc_p3 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qc_p3_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qc_p3_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qc_p3_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qc_p3_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qc_p3_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qc_p3_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qc_p3_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qc_p3_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qc_p3_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qc_p3_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qc_p3_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qb_p1 fifo_qd_p1 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qd_p1_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qd_p1_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qd_p1_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qd_p1_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qd_p1_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qd_p1_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qd_p1_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qd_p1_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qd_p1_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qd_p1_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qd_p1_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qb_p1 fifo_qd_p2 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qd_p2_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qd_p2_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qd_p2_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qd_p2_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qd_p2_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qd_p2_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qd_p2_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qd_p2_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qd_p2_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qd_p2_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qd_p2_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qb_p1 fifo_qd_p3 (
		.wrclock                          (pll_c0_clk),                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qd_p3_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qd_p3_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qd_p3_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qd_p3_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qd_p3_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qd_p3_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qd_p3_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qd_p3_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qd_p3_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qd_p3_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qd_p3_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_fifo_qb_p1 fifo_qe (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),            // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_qe_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_qe_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_qe_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_qe_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_qe_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_qe_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_qe_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_qe_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_qe_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_qe_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_qe_in_csr_readdata)   //         .readdata
	);

	FTOP_MSOC_jtag_uart_1a jtag_uart_1a (
		.clk            (pll_c0_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                      //               irq.irq
	);

	FTOP_MSOC_jtag_uart_1a jtag_uart_1f (
		.clk            (pll_c0_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver1_irq)                                  //               irq.irq
	);

	FTOP_MSOC_mem_info mem_info (
		.clk        (pll_c0_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_mem_info_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_mem_info_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_mem_info_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_mem_info_s1_write),      //       .write
		.readdata   (mm_interconnect_0_mem_info_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_mem_info_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_mem_info_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze     (1'b0)                                      // (terminated)
	);

	FTOP_MSOC_oc_ram_1f oc_ram_1f (
		.clk        (pll_c0_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_oc_ram_1f_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_oc_ram_1f_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_oc_ram_1f_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_oc_ram_1f_s1_write),      //       .write
		.readdata   (mm_interconnect_0_oc_ram_1f_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_oc_ram_1f_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_oc_ram_1f_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze     (1'b0)                                       // (terminated)
	);

	FTOP_MSOC_pll pll (
		.clk                (clk_clk),                                   //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),        // inclk_interface_reset.reset
		.read               (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0                 (pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                             //                    c1.clk
		.scandone           (),                                          //           (terminated)
		.scandataout        (),                                          //           (terminated)
		.phasecounterselect (4'b0000),                                   //           (terminated)
		.phaseupdown        (1'b0),                                      //           (terminated)
		.phasestep          (1'b0),                                      //           (terminated)
		.scanclk            (1'b0),                                      //           (terminated)
		.scanclkena         (1'b0),                                      //           (terminated)
		.scandata           (1'b0),                                      //           (terminated)
		.configupdate       (1'b0),                                      //           (terminated)
		.areset             (1'b0),                                      //           (terminated)
		.locked             (),                                          //           (terminated)
		.phasedone          ()                                           //           (terminated)
	);

	FTOP_MSOC_sdram_controller sdram_controller (
		.clk            (pll_c0_clk),                                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                           //      .export
	);

	FTOP_MSOC_sys_id_1a sys_id_1a (
		.clock    (pll_c0_clk),                                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                    //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_1a_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_1a_control_slave_address)   //              .address
	);

	FTOP_MSOC_sysid_1f sysid_1f (
		.clock    (pll_c0_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_1f_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_1f_control_slave_address)   //              .address
	);

	FTOP_MSOC_timer_1a timer_1a (
		.clk        (pll_c0_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_1a_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1a_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1a_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1a_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1a_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                  //   irq.irq
	);

	FTOP_MSOC_timer_1a timer_1f (
		.clk        (pll_c0_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_1f_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1f_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1f_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1f_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1f_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver0_irq)              //   irq.irq
	);

	FTOP_MSOC_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                         (clk_clk),                                                      //                                       clock_clk.clk
		.pll_c0_clk                                            (pll_c0_clk),                                                   //                                          pll_c0.clk
		.cpu_1a_reset_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                               //              cpu_1a_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                           // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_1a_data_master_address                            (cpu_1a_data_master_address),                                   //                              cpu_1a_data_master.address
		.cpu_1a_data_master_waitrequest                        (cpu_1a_data_master_waitrequest),                               //                                                .waitrequest
		.cpu_1a_data_master_byteenable                         (cpu_1a_data_master_byteenable),                                //                                                .byteenable
		.cpu_1a_data_master_read                               (cpu_1a_data_master_read),                                      //                                                .read
		.cpu_1a_data_master_readdata                           (cpu_1a_data_master_readdata),                                  //                                                .readdata
		.cpu_1a_data_master_write                              (cpu_1a_data_master_write),                                     //                                                .write
		.cpu_1a_data_master_writedata                          (cpu_1a_data_master_writedata),                                 //                                                .writedata
		.cpu_1a_data_master_debugaccess                        (cpu_1a_data_master_debugaccess),                               //                                                .debugaccess
		.cpu_1a_instruction_master_address                     (cpu_1a_instruction_master_address),                            //                       cpu_1a_instruction_master.address
		.cpu_1a_instruction_master_waitrequest                 (cpu_1a_instruction_master_waitrequest),                        //                                                .waitrequest
		.cpu_1a_instruction_master_read                        (cpu_1a_instruction_master_read),                               //                                                .read
		.cpu_1a_instruction_master_readdata                    (cpu_1a_instruction_master_readdata),                           //                                                .readdata
		.CPU_1b_p1_mm_bridge_0_m0_address                      (cpu_1b_p1_mm_bridge_0_m0_address),                             //                        CPU_1b_p1_mm_bridge_0_m0.address
		.CPU_1b_p1_mm_bridge_0_m0_waitrequest                  (cpu_1b_p1_mm_bridge_0_m0_waitrequest),                         //                                                .waitrequest
		.CPU_1b_p1_mm_bridge_0_m0_burstcount                   (cpu_1b_p1_mm_bridge_0_m0_burstcount),                          //                                                .burstcount
		.CPU_1b_p1_mm_bridge_0_m0_byteenable                   (cpu_1b_p1_mm_bridge_0_m0_byteenable),                          //                                                .byteenable
		.CPU_1b_p1_mm_bridge_0_m0_read                         (cpu_1b_p1_mm_bridge_0_m0_read),                                //                                                .read
		.CPU_1b_p1_mm_bridge_0_m0_readdata                     (cpu_1b_p1_mm_bridge_0_m0_readdata),                            //                                                .readdata
		.CPU_1b_p1_mm_bridge_0_m0_readdatavalid                (cpu_1b_p1_mm_bridge_0_m0_readdatavalid),                       //                                                .readdatavalid
		.CPU_1b_p1_mm_bridge_0_m0_write                        (cpu_1b_p1_mm_bridge_0_m0_write),                               //                                                .write
		.CPU_1b_p1_mm_bridge_0_m0_writedata                    (cpu_1b_p1_mm_bridge_0_m0_writedata),                           //                                                .writedata
		.CPU_1b_p1_mm_bridge_0_m0_debugaccess                  (cpu_1b_p1_mm_bridge_0_m0_debugaccess),                         //                                                .debugaccess
		.CPU_1b_p2_mm_bridge_0_m0_address                      (cpu_1b_p2_mm_bridge_0_m0_address),                             //                        CPU_1b_p2_mm_bridge_0_m0.address
		.CPU_1b_p2_mm_bridge_0_m0_waitrequest                  (cpu_1b_p2_mm_bridge_0_m0_waitrequest),                         //                                                .waitrequest
		.CPU_1b_p2_mm_bridge_0_m0_burstcount                   (cpu_1b_p2_mm_bridge_0_m0_burstcount),                          //                                                .burstcount
		.CPU_1b_p2_mm_bridge_0_m0_byteenable                   (cpu_1b_p2_mm_bridge_0_m0_byteenable),                          //                                                .byteenable
		.CPU_1b_p2_mm_bridge_0_m0_read                         (cpu_1b_p2_mm_bridge_0_m0_read),                                //                                                .read
		.CPU_1b_p2_mm_bridge_0_m0_readdata                     (cpu_1b_p2_mm_bridge_0_m0_readdata),                            //                                                .readdata
		.CPU_1b_p2_mm_bridge_0_m0_readdatavalid                (cpu_1b_p2_mm_bridge_0_m0_readdatavalid),                       //                                                .readdatavalid
		.CPU_1b_p2_mm_bridge_0_m0_write                        (cpu_1b_p2_mm_bridge_0_m0_write),                               //                                                .write
		.CPU_1b_p2_mm_bridge_0_m0_writedata                    (cpu_1b_p2_mm_bridge_0_m0_writedata),                           //                                                .writedata
		.CPU_1b_p2_mm_bridge_0_m0_debugaccess                  (cpu_1b_p2_mm_bridge_0_m0_debugaccess),                         //                                                .debugaccess
		.CPU_1b_p3_mm_bridge_0_m0_address                      (cpu_1b_p3_mm_bridge_0_m0_address),                             //                        CPU_1b_p3_mm_bridge_0_m0.address
		.CPU_1b_p3_mm_bridge_0_m0_waitrequest                  (cpu_1b_p3_mm_bridge_0_m0_waitrequest),                         //                                                .waitrequest
		.CPU_1b_p3_mm_bridge_0_m0_burstcount                   (cpu_1b_p3_mm_bridge_0_m0_burstcount),                          //                                                .burstcount
		.CPU_1b_p3_mm_bridge_0_m0_byteenable                   (cpu_1b_p3_mm_bridge_0_m0_byteenable),                          //                                                .byteenable
		.CPU_1b_p3_mm_bridge_0_m0_read                         (cpu_1b_p3_mm_bridge_0_m0_read),                                //                                                .read
		.CPU_1b_p3_mm_bridge_0_m0_readdata                     (cpu_1b_p3_mm_bridge_0_m0_readdata),                            //                                                .readdata
		.CPU_1b_p3_mm_bridge_0_m0_readdatavalid                (cpu_1b_p3_mm_bridge_0_m0_readdatavalid),                       //                                                .readdatavalid
		.CPU_1b_p3_mm_bridge_0_m0_write                        (cpu_1b_p3_mm_bridge_0_m0_write),                               //                                                .write
		.CPU_1b_p3_mm_bridge_0_m0_writedata                    (cpu_1b_p3_mm_bridge_0_m0_writedata),                           //                                                .writedata
		.CPU_1b_p3_mm_bridge_0_m0_debugaccess                  (cpu_1b_p3_mm_bridge_0_m0_debugaccess),                         //                                                .debugaccess
		.CPU_1c_p1_mm_bridge_0_m0_address                      (cpu_1c_p1_mm_bridge_0_m0_address),                             //                        CPU_1c_p1_mm_bridge_0_m0.address
		.CPU_1c_p1_mm_bridge_0_m0_waitrequest                  (cpu_1c_p1_mm_bridge_0_m0_waitrequest),                         //                                                .waitrequest
		.CPU_1c_p1_mm_bridge_0_m0_burstcount                   (cpu_1c_p1_mm_bridge_0_m0_burstcount),                          //                                                .burstcount
		.CPU_1c_p1_mm_bridge_0_m0_byteenable                   (cpu_1c_p1_mm_bridge_0_m0_byteenable),                          //                                                .byteenable
		.CPU_1c_p1_mm_bridge_0_m0_read                         (cpu_1c_p1_mm_bridge_0_m0_read),                                //                                                .read
		.CPU_1c_p1_mm_bridge_0_m0_readdata                     (cpu_1c_p1_mm_bridge_0_m0_readdata),                            //                                                .readdata
		.CPU_1c_p1_mm_bridge_0_m0_readdatavalid                (cpu_1c_p1_mm_bridge_0_m0_readdatavalid),                       //                                                .readdatavalid
		.CPU_1c_p1_mm_bridge_0_m0_write                        (cpu_1c_p1_mm_bridge_0_m0_write),                               //                                                .write
		.CPU_1c_p1_mm_bridge_0_m0_writedata                    (cpu_1c_p1_mm_bridge_0_m0_writedata),                           //                                                .writedata
		.CPU_1c_p1_mm_bridge_0_m0_debugaccess                  (cpu_1c_p1_mm_bridge_0_m0_debugaccess),                         //                                                .debugaccess
		.CPU_1c_p2_mm_bridge_0_m0_address                      (cpu_1c_p2_mm_bridge_0_m0_address),                             //                        CPU_1c_p2_mm_bridge_0_m0.address
		.CPU_1c_p2_mm_bridge_0_m0_waitrequest                  (cpu_1c_p2_mm_bridge_0_m0_waitrequest),                         //                                                .waitrequest
		.CPU_1c_p2_mm_bridge_0_m0_burstcount                   (cpu_1c_p2_mm_bridge_0_m0_burstcount),                          //                                                .burstcount
		.CPU_1c_p2_mm_bridge_0_m0_byteenable                   (cpu_1c_p2_mm_bridge_0_m0_byteenable),                          //                                                .byteenable
		.CPU_1c_p2_mm_bridge_0_m0_read                         (cpu_1c_p2_mm_bridge_0_m0_read),                                //                                                .read
		.CPU_1c_p2_mm_bridge_0_m0_readdata                     (cpu_1c_p2_mm_bridge_0_m0_readdata),                            //                                                .readdata
		.CPU_1c_p2_mm_bridge_0_m0_readdatavalid                (cpu_1c_p2_mm_bridge_0_m0_readdatavalid),                       //                                                .readdatavalid
		.CPU_1c_p2_mm_bridge_0_m0_write                        (cpu_1c_p2_mm_bridge_0_m0_write),                               //                                                .write
		.CPU_1c_p2_mm_bridge_0_m0_writedata                    (cpu_1c_p2_mm_bridge_0_m0_writedata),                           //                                                .writedata
		.CPU_1c_p2_mm_bridge_0_m0_debugaccess                  (cpu_1c_p2_mm_bridge_0_m0_debugaccess),                         //                                                .debugaccess
		.CPU_1c_p3_mm_bridge_0_m0_address                      (cpu_1c_p3_mm_bridge_0_m0_address),                             //                        CPU_1c_p3_mm_bridge_0_m0.address
		.CPU_1c_p3_mm_bridge_0_m0_waitrequest                  (cpu_1c_p3_mm_bridge_0_m0_waitrequest),                         //                                                .waitrequest
		.CPU_1c_p3_mm_bridge_0_m0_burstcount                   (cpu_1c_p3_mm_bridge_0_m0_burstcount),                          //                                                .burstcount
		.CPU_1c_p3_mm_bridge_0_m0_byteenable                   (cpu_1c_p3_mm_bridge_0_m0_byteenable),                          //                                                .byteenable
		.CPU_1c_p3_mm_bridge_0_m0_read                         (cpu_1c_p3_mm_bridge_0_m0_read),                                //                                                .read
		.CPU_1c_p3_mm_bridge_0_m0_readdata                     (cpu_1c_p3_mm_bridge_0_m0_readdata),                            //                                                .readdata
		.CPU_1c_p3_mm_bridge_0_m0_readdatavalid                (cpu_1c_p3_mm_bridge_0_m0_readdatavalid),                       //                                                .readdatavalid
		.CPU_1c_p3_mm_bridge_0_m0_write                        (cpu_1c_p3_mm_bridge_0_m0_write),                               //                                                .write
		.CPU_1c_p3_mm_bridge_0_m0_writedata                    (cpu_1c_p3_mm_bridge_0_m0_writedata),                           //                                                .writedata
		.CPU_1c_p3_mm_bridge_0_m0_debugaccess                  (cpu_1c_p3_mm_bridge_0_m0_debugaccess),                         //                                                .debugaccess
		.CPU_1d_p1_mm_bridge_0_m0_address                      (cpu_1d_p1_mm_bridge_0_m0_address),                             //                        CPU_1d_p1_mm_bridge_0_m0.address
		.CPU_1d_p1_mm_bridge_0_m0_waitrequest                  (cpu_1d_p1_mm_bridge_0_m0_waitrequest),                         //                                                .waitrequest
		.CPU_1d_p1_mm_bridge_0_m0_burstcount                   (cpu_1d_p1_mm_bridge_0_m0_burstcount),                          //                                                .burstcount
		.CPU_1d_p1_mm_bridge_0_m0_byteenable                   (cpu_1d_p1_mm_bridge_0_m0_byteenable),                          //                                                .byteenable
		.CPU_1d_p1_mm_bridge_0_m0_read                         (cpu_1d_p1_mm_bridge_0_m0_read),                                //                                                .read
		.CPU_1d_p1_mm_bridge_0_m0_readdata                     (cpu_1d_p1_mm_bridge_0_m0_readdata),                            //                                                .readdata
		.CPU_1d_p1_mm_bridge_0_m0_readdatavalid                (cpu_1d_p1_mm_bridge_0_m0_readdatavalid),                       //                                                .readdatavalid
		.CPU_1d_p1_mm_bridge_0_m0_write                        (cpu_1d_p1_mm_bridge_0_m0_write),                               //                                                .write
		.CPU_1d_p1_mm_bridge_0_m0_writedata                    (cpu_1d_p1_mm_bridge_0_m0_writedata),                           //                                                .writedata
		.CPU_1d_p1_mm_bridge_0_m0_debugaccess                  (cpu_1d_p1_mm_bridge_0_m0_debugaccess),                         //                                                .debugaccess
		.CPU_1d_p2_mm_bridge_0_m0_address                      (cpu_1d_p2_mm_bridge_0_m0_address),                             //                        CPU_1d_p2_mm_bridge_0_m0.address
		.CPU_1d_p2_mm_bridge_0_m0_waitrequest                  (cpu_1d_p2_mm_bridge_0_m0_waitrequest),                         //                                                .waitrequest
		.CPU_1d_p2_mm_bridge_0_m0_burstcount                   (cpu_1d_p2_mm_bridge_0_m0_burstcount),                          //                                                .burstcount
		.CPU_1d_p2_mm_bridge_0_m0_byteenable                   (cpu_1d_p2_mm_bridge_0_m0_byteenable),                          //                                                .byteenable
		.CPU_1d_p2_mm_bridge_0_m0_read                         (cpu_1d_p2_mm_bridge_0_m0_read),                                //                                                .read
		.CPU_1d_p2_mm_bridge_0_m0_readdata                     (cpu_1d_p2_mm_bridge_0_m0_readdata),                            //                                                .readdata
		.CPU_1d_p2_mm_bridge_0_m0_readdatavalid                (cpu_1d_p2_mm_bridge_0_m0_readdatavalid),                       //                                                .readdatavalid
		.CPU_1d_p2_mm_bridge_0_m0_write                        (cpu_1d_p2_mm_bridge_0_m0_write),                               //                                                .write
		.CPU_1d_p2_mm_bridge_0_m0_writedata                    (cpu_1d_p2_mm_bridge_0_m0_writedata),                           //                                                .writedata
		.CPU_1d_p2_mm_bridge_0_m0_debugaccess                  (cpu_1d_p2_mm_bridge_0_m0_debugaccess),                         //                                                .debugaccess
		.CPU_1d_p3_mm_bridge_0_m0_address                      (cpu_1d_p3_mm_bridge_0_m0_address),                             //                        CPU_1d_p3_mm_bridge_0_m0.address
		.CPU_1d_p3_mm_bridge_0_m0_waitrequest                  (cpu_1d_p3_mm_bridge_0_m0_waitrequest),                         //                                                .waitrequest
		.CPU_1d_p3_mm_bridge_0_m0_burstcount                   (cpu_1d_p3_mm_bridge_0_m0_burstcount),                          //                                                .burstcount
		.CPU_1d_p3_mm_bridge_0_m0_byteenable                   (cpu_1d_p3_mm_bridge_0_m0_byteenable),                          //                                                .byteenable
		.CPU_1d_p3_mm_bridge_0_m0_read                         (cpu_1d_p3_mm_bridge_0_m0_read),                                //                                                .read
		.CPU_1d_p3_mm_bridge_0_m0_readdata                     (cpu_1d_p3_mm_bridge_0_m0_readdata),                            //                                                .readdata
		.CPU_1d_p3_mm_bridge_0_m0_readdatavalid                (cpu_1d_p3_mm_bridge_0_m0_readdatavalid),                       //                                                .readdatavalid
		.CPU_1d_p3_mm_bridge_0_m0_write                        (cpu_1d_p3_mm_bridge_0_m0_write),                               //                                                .write
		.CPU_1d_p3_mm_bridge_0_m0_writedata                    (cpu_1d_p3_mm_bridge_0_m0_writedata),                           //                                                .writedata
		.CPU_1d_p3_mm_bridge_0_m0_debugaccess                  (cpu_1d_p3_mm_bridge_0_m0_debugaccess),                         //                                                .debugaccess
		.CPU_1e_mm_bridge_0_m0_address                         (cpu_1e_mm_bridge_0_m0_address),                                //                           CPU_1e_mm_bridge_0_m0.address
		.CPU_1e_mm_bridge_0_m0_waitrequest                     (cpu_1e_mm_bridge_0_m0_waitrequest),                            //                                                .waitrequest
		.CPU_1e_mm_bridge_0_m0_burstcount                      (cpu_1e_mm_bridge_0_m0_burstcount),                             //                                                .burstcount
		.CPU_1e_mm_bridge_0_m0_byteenable                      (cpu_1e_mm_bridge_0_m0_byteenable),                             //                                                .byteenable
		.CPU_1e_mm_bridge_0_m0_read                            (cpu_1e_mm_bridge_0_m0_read),                                   //                                                .read
		.CPU_1e_mm_bridge_0_m0_readdata                        (cpu_1e_mm_bridge_0_m0_readdata),                               //                                                .readdata
		.CPU_1e_mm_bridge_0_m0_readdatavalid                   (cpu_1e_mm_bridge_0_m0_readdatavalid),                          //                                                .readdatavalid
		.CPU_1e_mm_bridge_0_m0_write                           (cpu_1e_mm_bridge_0_m0_write),                                  //                                                .write
		.CPU_1e_mm_bridge_0_m0_writedata                       (cpu_1e_mm_bridge_0_m0_writedata),                              //                                                .writedata
		.CPU_1e_mm_bridge_0_m0_debugaccess                     (cpu_1e_mm_bridge_0_m0_debugaccess),                            //                                                .debugaccess
		.cpu_1f_data_master_address                            (cpu_1f_data_master_address),                                   //                              cpu_1f_data_master.address
		.cpu_1f_data_master_waitrequest                        (cpu_1f_data_master_waitrequest),                               //                                                .waitrequest
		.cpu_1f_data_master_byteenable                         (cpu_1f_data_master_byteenable),                                //                                                .byteenable
		.cpu_1f_data_master_read                               (cpu_1f_data_master_read),                                      //                                                .read
		.cpu_1f_data_master_readdata                           (cpu_1f_data_master_readdata),                                  //                                                .readdata
		.cpu_1f_data_master_write                              (cpu_1f_data_master_write),                                     //                                                .write
		.cpu_1f_data_master_writedata                          (cpu_1f_data_master_writedata),                                 //                                                .writedata
		.cpu_1f_data_master_debugaccess                        (cpu_1f_data_master_debugaccess),                               //                                                .debugaccess
		.cpu_1f_instruction_master_address                     (cpu_1f_instruction_master_address),                            //                       cpu_1f_instruction_master.address
		.cpu_1f_instruction_master_waitrequest                 (cpu_1f_instruction_master_waitrequest),                        //                                                .waitrequest
		.cpu_1f_instruction_master_read                        (cpu_1f_instruction_master_read),                               //                                                .read
		.cpu_1f_instruction_master_readdata                    (cpu_1f_instruction_master_readdata),                           //                                                .readdata
		.cpu_1a_debug_mem_slave_address                        (mm_interconnect_0_cpu_1a_debug_mem_slave_address),             //                          cpu_1a_debug_mem_slave.address
		.cpu_1a_debug_mem_slave_write                          (mm_interconnect_0_cpu_1a_debug_mem_slave_write),               //                                                .write
		.cpu_1a_debug_mem_slave_read                           (mm_interconnect_0_cpu_1a_debug_mem_slave_read),                //                                                .read
		.cpu_1a_debug_mem_slave_readdata                       (mm_interconnect_0_cpu_1a_debug_mem_slave_readdata),            //                                                .readdata
		.cpu_1a_debug_mem_slave_writedata                      (mm_interconnect_0_cpu_1a_debug_mem_slave_writedata),           //                                                .writedata
		.cpu_1a_debug_mem_slave_byteenable                     (mm_interconnect_0_cpu_1a_debug_mem_slave_byteenable),          //                                                .byteenable
		.cpu_1a_debug_mem_slave_waitrequest                    (mm_interconnect_0_cpu_1a_debug_mem_slave_waitrequest),         //                                                .waitrequest
		.cpu_1a_debug_mem_slave_debugaccess                    (mm_interconnect_0_cpu_1a_debug_mem_slave_debugaccess),         //                                                .debugaccess
		.cpu_1f_debug_mem_slave_address                        (mm_interconnect_0_cpu_1f_debug_mem_slave_address),             //                          cpu_1f_debug_mem_slave.address
		.cpu_1f_debug_mem_slave_write                          (mm_interconnect_0_cpu_1f_debug_mem_slave_write),               //                                                .write
		.cpu_1f_debug_mem_slave_read                           (mm_interconnect_0_cpu_1f_debug_mem_slave_read),                //                                                .read
		.cpu_1f_debug_mem_slave_readdata                       (mm_interconnect_0_cpu_1f_debug_mem_slave_readdata),            //                                                .readdata
		.cpu_1f_debug_mem_slave_writedata                      (mm_interconnect_0_cpu_1f_debug_mem_slave_writedata),           //                                                .writedata
		.cpu_1f_debug_mem_slave_byteenable                     (mm_interconnect_0_cpu_1f_debug_mem_slave_byteenable),          //                                                .byteenable
		.cpu_1f_debug_mem_slave_waitrequest                    (mm_interconnect_0_cpu_1f_debug_mem_slave_waitrequest),         //                                                .waitrequest
		.cpu_1f_debug_mem_slave_debugaccess                    (mm_interconnect_0_cpu_1f_debug_mem_slave_debugaccess),         //                                                .debugaccess
		.fifo_qa_p1_in_write                                   (mm_interconnect_0_fifo_qa_p1_in_write),                        //                                   fifo_qa_p1_in.write
		.fifo_qa_p1_in_writedata                               (mm_interconnect_0_fifo_qa_p1_in_writedata),                    //                                                .writedata
		.fifo_qa_p1_in_waitrequest                             (mm_interconnect_0_fifo_qa_p1_in_waitrequest),                  //                                                .waitrequest
		.fifo_qa_p1_in_csr_address                             (mm_interconnect_0_fifo_qa_p1_in_csr_address),                  //                               fifo_qa_p1_in_csr.address
		.fifo_qa_p1_in_csr_write                               (mm_interconnect_0_fifo_qa_p1_in_csr_write),                    //                                                .write
		.fifo_qa_p1_in_csr_read                                (mm_interconnect_0_fifo_qa_p1_in_csr_read),                     //                                                .read
		.fifo_qa_p1_in_csr_readdata                            (mm_interconnect_0_fifo_qa_p1_in_csr_readdata),                 //                                                .readdata
		.fifo_qa_p1_in_csr_writedata                           (mm_interconnect_0_fifo_qa_p1_in_csr_writedata),                //                                                .writedata
		.fifo_qa_p1_out_read                                   (mm_interconnect_0_fifo_qa_p1_out_read),                        //                                  fifo_qa_p1_out.read
		.fifo_qa_p1_out_readdata                               (mm_interconnect_0_fifo_qa_p1_out_readdata),                    //                                                .readdata
		.fifo_qa_p1_out_waitrequest                            (mm_interconnect_0_fifo_qa_p1_out_waitrequest),                 //                                                .waitrequest
		.fifo_qa_p2_in_write                                   (mm_interconnect_0_fifo_qa_p2_in_write),                        //                                   fifo_qa_p2_in.write
		.fifo_qa_p2_in_writedata                               (mm_interconnect_0_fifo_qa_p2_in_writedata),                    //                                                .writedata
		.fifo_qa_p2_in_waitrequest                             (mm_interconnect_0_fifo_qa_p2_in_waitrequest),                  //                                                .waitrequest
		.fifo_qa_p2_in_csr_address                             (mm_interconnect_0_fifo_qa_p2_in_csr_address),                  //                               fifo_qa_p2_in_csr.address
		.fifo_qa_p2_in_csr_write                               (mm_interconnect_0_fifo_qa_p2_in_csr_write),                    //                                                .write
		.fifo_qa_p2_in_csr_read                                (mm_interconnect_0_fifo_qa_p2_in_csr_read),                     //                                                .read
		.fifo_qa_p2_in_csr_readdata                            (mm_interconnect_0_fifo_qa_p2_in_csr_readdata),                 //                                                .readdata
		.fifo_qa_p2_in_csr_writedata                           (mm_interconnect_0_fifo_qa_p2_in_csr_writedata),                //                                                .writedata
		.fifo_qa_p2_out_read                                   (mm_interconnect_0_fifo_qa_p2_out_read),                        //                                  fifo_qa_p2_out.read
		.fifo_qa_p2_out_readdata                               (mm_interconnect_0_fifo_qa_p2_out_readdata),                    //                                                .readdata
		.fifo_qa_p2_out_waitrequest                            (mm_interconnect_0_fifo_qa_p2_out_waitrequest),                 //                                                .waitrequest
		.fifo_qa_p3_in_write                                   (mm_interconnect_0_fifo_qa_p3_in_write),                        //                                   fifo_qa_p3_in.write
		.fifo_qa_p3_in_writedata                               (mm_interconnect_0_fifo_qa_p3_in_writedata),                    //                                                .writedata
		.fifo_qa_p3_in_waitrequest                             (mm_interconnect_0_fifo_qa_p3_in_waitrequest),                  //                                                .waitrequest
		.fifo_qa_p3_in_csr_address                             (mm_interconnect_0_fifo_qa_p3_in_csr_address),                  //                               fifo_qa_p3_in_csr.address
		.fifo_qa_p3_in_csr_write                               (mm_interconnect_0_fifo_qa_p3_in_csr_write),                    //                                                .write
		.fifo_qa_p3_in_csr_read                                (mm_interconnect_0_fifo_qa_p3_in_csr_read),                     //                                                .read
		.fifo_qa_p3_in_csr_readdata                            (mm_interconnect_0_fifo_qa_p3_in_csr_readdata),                 //                                                .readdata
		.fifo_qa_p3_in_csr_writedata                           (mm_interconnect_0_fifo_qa_p3_in_csr_writedata),                //                                                .writedata
		.fifo_qa_p3_out_read                                   (mm_interconnect_0_fifo_qa_p3_out_read),                        //                                  fifo_qa_p3_out.read
		.fifo_qa_p3_out_readdata                               (mm_interconnect_0_fifo_qa_p3_out_readdata),                    //                                                .readdata
		.fifo_qa_p3_out_waitrequest                            (mm_interconnect_0_fifo_qa_p3_out_waitrequest),                 //                                                .waitrequest
		.fifo_qb_p1_in_write                                   (mm_interconnect_0_fifo_qb_p1_in_write),                        //                                   fifo_qb_p1_in.write
		.fifo_qb_p1_in_writedata                               (mm_interconnect_0_fifo_qb_p1_in_writedata),                    //                                                .writedata
		.fifo_qb_p1_in_waitrequest                             (mm_interconnect_0_fifo_qb_p1_in_waitrequest),                  //                                                .waitrequest
		.fifo_qb_p1_in_csr_address                             (mm_interconnect_0_fifo_qb_p1_in_csr_address),                  //                               fifo_qb_p1_in_csr.address
		.fifo_qb_p1_in_csr_write                               (mm_interconnect_0_fifo_qb_p1_in_csr_write),                    //                                                .write
		.fifo_qb_p1_in_csr_read                                (mm_interconnect_0_fifo_qb_p1_in_csr_read),                     //                                                .read
		.fifo_qb_p1_in_csr_readdata                            (mm_interconnect_0_fifo_qb_p1_in_csr_readdata),                 //                                                .readdata
		.fifo_qb_p1_in_csr_writedata                           (mm_interconnect_0_fifo_qb_p1_in_csr_writedata),                //                                                .writedata
		.fifo_qb_p1_out_read                                   (mm_interconnect_0_fifo_qb_p1_out_read),                        //                                  fifo_qb_p1_out.read
		.fifo_qb_p1_out_readdata                               (mm_interconnect_0_fifo_qb_p1_out_readdata),                    //                                                .readdata
		.fifo_qb_p1_out_waitrequest                            (mm_interconnect_0_fifo_qb_p1_out_waitrequest),                 //                                                .waitrequest
		.fifo_qb_p2_in_write                                   (mm_interconnect_0_fifo_qb_p2_in_write),                        //                                   fifo_qb_p2_in.write
		.fifo_qb_p2_in_writedata                               (mm_interconnect_0_fifo_qb_p2_in_writedata),                    //                                                .writedata
		.fifo_qb_p2_in_waitrequest                             (mm_interconnect_0_fifo_qb_p2_in_waitrequest),                  //                                                .waitrequest
		.fifo_qb_p2_in_csr_address                             (mm_interconnect_0_fifo_qb_p2_in_csr_address),                  //                               fifo_qb_p2_in_csr.address
		.fifo_qb_p2_in_csr_write                               (mm_interconnect_0_fifo_qb_p2_in_csr_write),                    //                                                .write
		.fifo_qb_p2_in_csr_read                                (mm_interconnect_0_fifo_qb_p2_in_csr_read),                     //                                                .read
		.fifo_qb_p2_in_csr_readdata                            (mm_interconnect_0_fifo_qb_p2_in_csr_readdata),                 //                                                .readdata
		.fifo_qb_p2_in_csr_writedata                           (mm_interconnect_0_fifo_qb_p2_in_csr_writedata),                //                                                .writedata
		.fifo_qb_p2_out_read                                   (mm_interconnect_0_fifo_qb_p2_out_read),                        //                                  fifo_qb_p2_out.read
		.fifo_qb_p2_out_readdata                               (mm_interconnect_0_fifo_qb_p2_out_readdata),                    //                                                .readdata
		.fifo_qb_p2_out_waitrequest                            (mm_interconnect_0_fifo_qb_p2_out_waitrequest),                 //                                                .waitrequest
		.fifo_qb_p3_in_write                                   (mm_interconnect_0_fifo_qb_p3_in_write),                        //                                   fifo_qb_p3_in.write
		.fifo_qb_p3_in_writedata                               (mm_interconnect_0_fifo_qb_p3_in_writedata),                    //                                                .writedata
		.fifo_qb_p3_in_waitrequest                             (mm_interconnect_0_fifo_qb_p3_in_waitrequest),                  //                                                .waitrequest
		.fifo_qb_p3_in_csr_address                             (mm_interconnect_0_fifo_qb_p3_in_csr_address),                  //                               fifo_qb_p3_in_csr.address
		.fifo_qb_p3_in_csr_write                               (mm_interconnect_0_fifo_qb_p3_in_csr_write),                    //                                                .write
		.fifo_qb_p3_in_csr_read                                (mm_interconnect_0_fifo_qb_p3_in_csr_read),                     //                                                .read
		.fifo_qb_p3_in_csr_readdata                            (mm_interconnect_0_fifo_qb_p3_in_csr_readdata),                 //                                                .readdata
		.fifo_qb_p3_in_csr_writedata                           (mm_interconnect_0_fifo_qb_p3_in_csr_writedata),                //                                                .writedata
		.fifo_qb_p3_out_read                                   (mm_interconnect_0_fifo_qb_p3_out_read),                        //                                  fifo_qb_p3_out.read
		.fifo_qb_p3_out_readdata                               (mm_interconnect_0_fifo_qb_p3_out_readdata),                    //                                                .readdata
		.fifo_qb_p3_out_waitrequest                            (mm_interconnect_0_fifo_qb_p3_out_waitrequest),                 //                                                .waitrequest
		.fifo_qc_p1_in_write                                   (mm_interconnect_0_fifo_qc_p1_in_write),                        //                                   fifo_qc_p1_in.write
		.fifo_qc_p1_in_writedata                               (mm_interconnect_0_fifo_qc_p1_in_writedata),                    //                                                .writedata
		.fifo_qc_p1_in_waitrequest                             (mm_interconnect_0_fifo_qc_p1_in_waitrequest),                  //                                                .waitrequest
		.fifo_qc_p1_in_csr_address                             (mm_interconnect_0_fifo_qc_p1_in_csr_address),                  //                               fifo_qc_p1_in_csr.address
		.fifo_qc_p1_in_csr_write                               (mm_interconnect_0_fifo_qc_p1_in_csr_write),                    //                                                .write
		.fifo_qc_p1_in_csr_read                                (mm_interconnect_0_fifo_qc_p1_in_csr_read),                     //                                                .read
		.fifo_qc_p1_in_csr_readdata                            (mm_interconnect_0_fifo_qc_p1_in_csr_readdata),                 //                                                .readdata
		.fifo_qc_p1_in_csr_writedata                           (mm_interconnect_0_fifo_qc_p1_in_csr_writedata),                //                                                .writedata
		.fifo_qc_p1_out_read                                   (mm_interconnect_0_fifo_qc_p1_out_read),                        //                                  fifo_qc_p1_out.read
		.fifo_qc_p1_out_readdata                               (mm_interconnect_0_fifo_qc_p1_out_readdata),                    //                                                .readdata
		.fifo_qc_p1_out_waitrequest                            (mm_interconnect_0_fifo_qc_p1_out_waitrequest),                 //                                                .waitrequest
		.fifo_qc_p2_in_write                                   (mm_interconnect_0_fifo_qc_p2_in_write),                        //                                   fifo_qc_p2_in.write
		.fifo_qc_p2_in_writedata                               (mm_interconnect_0_fifo_qc_p2_in_writedata),                    //                                                .writedata
		.fifo_qc_p2_in_waitrequest                             (mm_interconnect_0_fifo_qc_p2_in_waitrequest),                  //                                                .waitrequest
		.fifo_qc_p2_in_csr_address                             (mm_interconnect_0_fifo_qc_p2_in_csr_address),                  //                               fifo_qc_p2_in_csr.address
		.fifo_qc_p2_in_csr_write                               (mm_interconnect_0_fifo_qc_p2_in_csr_write),                    //                                                .write
		.fifo_qc_p2_in_csr_read                                (mm_interconnect_0_fifo_qc_p2_in_csr_read),                     //                                                .read
		.fifo_qc_p2_in_csr_readdata                            (mm_interconnect_0_fifo_qc_p2_in_csr_readdata),                 //                                                .readdata
		.fifo_qc_p2_in_csr_writedata                           (mm_interconnect_0_fifo_qc_p2_in_csr_writedata),                //                                                .writedata
		.fifo_qc_p2_out_read                                   (mm_interconnect_0_fifo_qc_p2_out_read),                        //                                  fifo_qc_p2_out.read
		.fifo_qc_p2_out_readdata                               (mm_interconnect_0_fifo_qc_p2_out_readdata),                    //                                                .readdata
		.fifo_qc_p2_out_waitrequest                            (mm_interconnect_0_fifo_qc_p2_out_waitrequest),                 //                                                .waitrequest
		.fifo_qc_p3_in_write                                   (mm_interconnect_0_fifo_qc_p3_in_write),                        //                                   fifo_qc_p3_in.write
		.fifo_qc_p3_in_writedata                               (mm_interconnect_0_fifo_qc_p3_in_writedata),                    //                                                .writedata
		.fifo_qc_p3_in_waitrequest                             (mm_interconnect_0_fifo_qc_p3_in_waitrequest),                  //                                                .waitrequest
		.fifo_qc_p3_in_csr_address                             (mm_interconnect_0_fifo_qc_p3_in_csr_address),                  //                               fifo_qc_p3_in_csr.address
		.fifo_qc_p3_in_csr_write                               (mm_interconnect_0_fifo_qc_p3_in_csr_write),                    //                                                .write
		.fifo_qc_p3_in_csr_read                                (mm_interconnect_0_fifo_qc_p3_in_csr_read),                     //                                                .read
		.fifo_qc_p3_in_csr_readdata                            (mm_interconnect_0_fifo_qc_p3_in_csr_readdata),                 //                                                .readdata
		.fifo_qc_p3_in_csr_writedata                           (mm_interconnect_0_fifo_qc_p3_in_csr_writedata),                //                                                .writedata
		.fifo_qc_p3_out_read                                   (mm_interconnect_0_fifo_qc_p3_out_read),                        //                                  fifo_qc_p3_out.read
		.fifo_qc_p3_out_readdata                               (mm_interconnect_0_fifo_qc_p3_out_readdata),                    //                                                .readdata
		.fifo_qc_p3_out_waitrequest                            (mm_interconnect_0_fifo_qc_p3_out_waitrequest),                 //                                                .waitrequest
		.fifo_qd_p1_in_write                                   (mm_interconnect_0_fifo_qd_p1_in_write),                        //                                   fifo_qd_p1_in.write
		.fifo_qd_p1_in_writedata                               (mm_interconnect_0_fifo_qd_p1_in_writedata),                    //                                                .writedata
		.fifo_qd_p1_in_waitrequest                             (mm_interconnect_0_fifo_qd_p1_in_waitrequest),                  //                                                .waitrequest
		.fifo_qd_p1_in_csr_address                             (mm_interconnect_0_fifo_qd_p1_in_csr_address),                  //                               fifo_qd_p1_in_csr.address
		.fifo_qd_p1_in_csr_write                               (mm_interconnect_0_fifo_qd_p1_in_csr_write),                    //                                                .write
		.fifo_qd_p1_in_csr_read                                (mm_interconnect_0_fifo_qd_p1_in_csr_read),                     //                                                .read
		.fifo_qd_p1_in_csr_readdata                            (mm_interconnect_0_fifo_qd_p1_in_csr_readdata),                 //                                                .readdata
		.fifo_qd_p1_in_csr_writedata                           (mm_interconnect_0_fifo_qd_p1_in_csr_writedata),                //                                                .writedata
		.fifo_qd_p1_out_read                                   (mm_interconnect_0_fifo_qd_p1_out_read),                        //                                  fifo_qd_p1_out.read
		.fifo_qd_p1_out_readdata                               (mm_interconnect_0_fifo_qd_p1_out_readdata),                    //                                                .readdata
		.fifo_qd_p1_out_waitrequest                            (mm_interconnect_0_fifo_qd_p1_out_waitrequest),                 //                                                .waitrequest
		.fifo_qd_p2_in_write                                   (mm_interconnect_0_fifo_qd_p2_in_write),                        //                                   fifo_qd_p2_in.write
		.fifo_qd_p2_in_writedata                               (mm_interconnect_0_fifo_qd_p2_in_writedata),                    //                                                .writedata
		.fifo_qd_p2_in_waitrequest                             (mm_interconnect_0_fifo_qd_p2_in_waitrequest),                  //                                                .waitrequest
		.fifo_qd_p2_in_csr_address                             (mm_interconnect_0_fifo_qd_p2_in_csr_address),                  //                               fifo_qd_p2_in_csr.address
		.fifo_qd_p2_in_csr_write                               (mm_interconnect_0_fifo_qd_p2_in_csr_write),                    //                                                .write
		.fifo_qd_p2_in_csr_read                                (mm_interconnect_0_fifo_qd_p2_in_csr_read),                     //                                                .read
		.fifo_qd_p2_in_csr_readdata                            (mm_interconnect_0_fifo_qd_p2_in_csr_readdata),                 //                                                .readdata
		.fifo_qd_p2_in_csr_writedata                           (mm_interconnect_0_fifo_qd_p2_in_csr_writedata),                //                                                .writedata
		.fifo_qd_p2_out_read                                   (mm_interconnect_0_fifo_qd_p2_out_read),                        //                                  fifo_qd_p2_out.read
		.fifo_qd_p2_out_readdata                               (mm_interconnect_0_fifo_qd_p2_out_readdata),                    //                                                .readdata
		.fifo_qd_p2_out_waitrequest                            (mm_interconnect_0_fifo_qd_p2_out_waitrequest),                 //                                                .waitrequest
		.fifo_qd_p3_in_write                                   (mm_interconnect_0_fifo_qd_p3_in_write),                        //                                   fifo_qd_p3_in.write
		.fifo_qd_p3_in_writedata                               (mm_interconnect_0_fifo_qd_p3_in_writedata),                    //                                                .writedata
		.fifo_qd_p3_in_waitrequest                             (mm_interconnect_0_fifo_qd_p3_in_waitrequest),                  //                                                .waitrequest
		.fifo_qd_p3_in_csr_address                             (mm_interconnect_0_fifo_qd_p3_in_csr_address),                  //                               fifo_qd_p3_in_csr.address
		.fifo_qd_p3_in_csr_write                               (mm_interconnect_0_fifo_qd_p3_in_csr_write),                    //                                                .write
		.fifo_qd_p3_in_csr_read                                (mm_interconnect_0_fifo_qd_p3_in_csr_read),                     //                                                .read
		.fifo_qd_p3_in_csr_readdata                            (mm_interconnect_0_fifo_qd_p3_in_csr_readdata),                 //                                                .readdata
		.fifo_qd_p3_in_csr_writedata                           (mm_interconnect_0_fifo_qd_p3_in_csr_writedata),                //                                                .writedata
		.fifo_qd_p3_out_read                                   (mm_interconnect_0_fifo_qd_p3_out_read),                        //                                  fifo_qd_p3_out.read
		.fifo_qd_p3_out_readdata                               (mm_interconnect_0_fifo_qd_p3_out_readdata),                    //                                                .readdata
		.fifo_qd_p3_out_waitrequest                            (mm_interconnect_0_fifo_qd_p3_out_waitrequest),                 //                                                .waitrequest
		.fifo_qe_in_write                                      (mm_interconnect_0_fifo_qe_in_write),                           //                                      fifo_qe_in.write
		.fifo_qe_in_writedata                                  (mm_interconnect_0_fifo_qe_in_writedata),                       //                                                .writedata
		.fifo_qe_in_waitrequest                                (mm_interconnect_0_fifo_qe_in_waitrequest),                     //                                                .waitrequest
		.fifo_qe_in_csr_address                                (mm_interconnect_0_fifo_qe_in_csr_address),                     //                                  fifo_qe_in_csr.address
		.fifo_qe_in_csr_write                                  (mm_interconnect_0_fifo_qe_in_csr_write),                       //                                                .write
		.fifo_qe_in_csr_read                                   (mm_interconnect_0_fifo_qe_in_csr_read),                        //                                                .read
		.fifo_qe_in_csr_readdata                               (mm_interconnect_0_fifo_qe_in_csr_readdata),                    //                                                .readdata
		.fifo_qe_in_csr_writedata                              (mm_interconnect_0_fifo_qe_in_csr_writedata),                   //                                                .writedata
		.fifo_qe_out_read                                      (mm_interconnect_0_fifo_qe_out_read),                           //                                     fifo_qe_out.read
		.fifo_qe_out_readdata                                  (mm_interconnect_0_fifo_qe_out_readdata),                       //                                                .readdata
		.fifo_qe_out_waitrequest                               (mm_interconnect_0_fifo_qe_out_waitrequest),                    //                                                .waitrequest
		.jtag_uart_1a_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_address),     //                  jtag_uart_1a_avalon_jtag_slave.address
		.jtag_uart_1a_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_1a_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_1a_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_1a_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_1a_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_1a_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_1a_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.jtag_uart_1f_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_address),     //                  jtag_uart_1f_avalon_jtag_slave.address
		.jtag_uart_1f_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_1f_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_1f_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_1f_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_1f_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_1f_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.mem_info_s1_address                                   (mm_interconnect_0_mem_info_s1_address),                        //                                     mem_info_s1.address
		.mem_info_s1_write                                     (mm_interconnect_0_mem_info_s1_write),                          //                                                .write
		.mem_info_s1_readdata                                  (mm_interconnect_0_mem_info_s1_readdata),                       //                                                .readdata
		.mem_info_s1_writedata                                 (mm_interconnect_0_mem_info_s1_writedata),                      //                                                .writedata
		.mem_info_s1_byteenable                                (mm_interconnect_0_mem_info_s1_byteenable),                     //                                                .byteenable
		.mem_info_s1_chipselect                                (mm_interconnect_0_mem_info_s1_chipselect),                     //                                                .chipselect
		.mem_info_s1_clken                                     (mm_interconnect_0_mem_info_s1_clken),                          //                                                .clken
		.oc_ram_1f_s1_address                                  (mm_interconnect_0_oc_ram_1f_s1_address),                       //                                    oc_ram_1f_s1.address
		.oc_ram_1f_s1_write                                    (mm_interconnect_0_oc_ram_1f_s1_write),                         //                                                .write
		.oc_ram_1f_s1_readdata                                 (mm_interconnect_0_oc_ram_1f_s1_readdata),                      //                                                .readdata
		.oc_ram_1f_s1_writedata                                (mm_interconnect_0_oc_ram_1f_s1_writedata),                     //                                                .writedata
		.oc_ram_1f_s1_byteenable                               (mm_interconnect_0_oc_ram_1f_s1_byteenable),                    //                                                .byteenable
		.oc_ram_1f_s1_chipselect                               (mm_interconnect_0_oc_ram_1f_s1_chipselect),                    //                                                .chipselect
		.oc_ram_1f_s1_clken                                    (mm_interconnect_0_oc_ram_1f_s1_clken),                         //                                                .clken
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                      //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                        //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                         //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                     //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                    //                                                .writedata
		.sdram_controller_s1_address                           (mm_interconnect_0_sdram_controller_s1_address),                //                             sdram_controller_s1.address
		.sdram_controller_s1_write                             (mm_interconnect_0_sdram_controller_s1_write),                  //                                                .write
		.sdram_controller_s1_read                              (mm_interconnect_0_sdram_controller_s1_read),                   //                                                .read
		.sdram_controller_s1_readdata                          (mm_interconnect_0_sdram_controller_s1_readdata),               //                                                .readdata
		.sdram_controller_s1_writedata                         (mm_interconnect_0_sdram_controller_s1_writedata),              //                                                .writedata
		.sdram_controller_s1_byteenable                        (mm_interconnect_0_sdram_controller_s1_byteenable),             //                                                .byteenable
		.sdram_controller_s1_readdatavalid                     (mm_interconnect_0_sdram_controller_s1_readdatavalid),          //                                                .readdatavalid
		.sdram_controller_s1_waitrequest                       (mm_interconnect_0_sdram_controller_s1_waitrequest),            //                                                .waitrequest
		.sdram_controller_s1_chipselect                        (mm_interconnect_0_sdram_controller_s1_chipselect),             //                                                .chipselect
		.sys_id_1a_control_slave_address                       (mm_interconnect_0_sys_id_1a_control_slave_address),            //                         sys_id_1a_control_slave.address
		.sys_id_1a_control_slave_readdata                      (mm_interconnect_0_sys_id_1a_control_slave_readdata),           //                                                .readdata
		.sysid_1f_control_slave_address                        (mm_interconnect_0_sysid_1f_control_slave_address),             //                          sysid_1f_control_slave.address
		.sysid_1f_control_slave_readdata                       (mm_interconnect_0_sysid_1f_control_slave_readdata),            //                                                .readdata
		.timer_1a_s1_address                                   (mm_interconnect_0_timer_1a_s1_address),                        //                                     timer_1a_s1.address
		.timer_1a_s1_write                                     (mm_interconnect_0_timer_1a_s1_write),                          //                                                .write
		.timer_1a_s1_readdata                                  (mm_interconnect_0_timer_1a_s1_readdata),                       //                                                .readdata
		.timer_1a_s1_writedata                                 (mm_interconnect_0_timer_1a_s1_writedata),                      //                                                .writedata
		.timer_1a_s1_chipselect                                (mm_interconnect_0_timer_1a_s1_chipselect),                     //                                                .chipselect
		.timer_1f_s1_address                                   (mm_interconnect_0_timer_1f_s1_address),                        //                                     timer_1f_s1.address
		.timer_1f_s1_write                                     (mm_interconnect_0_timer_1f_s1_write),                          //                                                .write
		.timer_1f_s1_readdata                                  (mm_interconnect_0_timer_1f_s1_readdata),                       //                                                .readdata
		.timer_1f_s1_writedata                                 (mm_interconnect_0_timer_1f_s1_writedata),                      //                                                .writedata
		.timer_1f_s1_chipselect                                (mm_interconnect_0_timer_1f_s1_chipselect)                      //                                                .chipselect
	);

	FTOP_MSOC_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_1a_irq_irq)                  //    sender.irq
	);

	FTOP_MSOC_irq_mapper irq_mapper_001 (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),   // receiver1.irq
		.sender_irq    (cpu_1f_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_1a_debug_reset_request_reset),   // reset_in1.reset
		.reset_in2      (cpu_1f_debug_reset_request_reset),   // reset_in2.reset
		.clk            (pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_1a_debug_reset_request_reset),   // reset_in1.reset
		.reset_in2      (cpu_1f_debug_reset_request_reset),   // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
