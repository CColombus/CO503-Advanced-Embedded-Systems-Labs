// TOP_MSOC.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module TOP_MSOC (
		input  wire        clk_clk,                     //                   clk.clk
		input  wire        reset_reset_n,               //                 reset.reset_n
		output wire        sdram_clk_clk,               //             sdram_clk.clk
		output wire [12:0] sdram_controller_wire_addr,  // sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,    //                      .ba
		output wire        sdram_controller_wire_cas_n, //                      .cas_n
		output wire        sdram_controller_wire_cke,   //                      .cke
		output wire        sdram_controller_wire_cs_n,  //                      .cs_n
		inout  wire [31:0] sdram_controller_wire_dq,    //                      .dq
		output wire [3:0]  sdram_controller_wire_dqm,   //                      .dqm
		output wire        sdram_controller_wire_ras_n, //                      .ras_n
		output wire        sdram_controller_wire_we_n   //                      .we_n
	);

	wire         pll_c0_clk;                                                   // pll:c0 -> [CPU_1b:clock_bridge_0_in_clk_clk, CPU_1c:clock_bridge_0_in_clk_clk, CPU_1d:clock_bridge_0_in_clk_clk, CPU_1e:clock_bridge_0_in_clk_clk, cpu:clk, cpu_1f:clk, fifo_1b:wrclock, fifo_1c:wrclock, fifo_1d:wrclock, fifo_1e:wrclock, fifo_q_1:wrclock, fifo_q_2:wrclock, fifo_q_3:wrclock, fifo_q_4:wrclock, fifo_q_5:wrclock, fifo_q_6:wrclock, irq_mapper:clk, irq_mapper_001:clk, jtag_uart:clk, jtag_uart_1f:clk, mm_interconnect_0:pll_c0_clk, rst_controller:clk, rst_controller_001:clk, sdram_controller:clk, sys_id:clock, sysid_1f:clock, timer:clk, timer_1f:clk]
	wire  [31:0] cpu_data_master_readdata;                                     // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                  // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                  // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                      // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                   // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                         // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                        // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                    // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_1f_data_master_readdata;                                  // mm_interconnect_0:cpu_1f_data_master_readdata -> cpu_1f:d_readdata
	wire         cpu_1f_data_master_waitrequest;                               // mm_interconnect_0:cpu_1f_data_master_waitrequest -> cpu_1f:d_waitrequest
	wire         cpu_1f_data_master_debugaccess;                               // cpu_1f:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1f_data_master_debugaccess
	wire  [27:0] cpu_1f_data_master_address;                                   // cpu_1f:d_address -> mm_interconnect_0:cpu_1f_data_master_address
	wire   [3:0] cpu_1f_data_master_byteenable;                                // cpu_1f:d_byteenable -> mm_interconnect_0:cpu_1f_data_master_byteenable
	wire         cpu_1f_data_master_read;                                      // cpu_1f:d_read -> mm_interconnect_0:cpu_1f_data_master_read
	wire         cpu_1f_data_master_write;                                     // cpu_1f:d_write -> mm_interconnect_0:cpu_1f_data_master_write
	wire  [31:0] cpu_1f_data_master_writedata;                                 // cpu_1f:d_writedata -> mm_interconnect_0:cpu_1f_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                              // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                           // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                               // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                  // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_1f_instruction_master_readdata;                           // mm_interconnect_0:cpu_1f_instruction_master_readdata -> cpu_1f:i_readdata
	wire         cpu_1f_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_1f_instruction_master_waitrequest -> cpu_1f:i_waitrequest
	wire  [27:0] cpu_1f_instruction_master_address;                            // cpu_1f:i_address -> mm_interconnect_0:cpu_1f_instruction_master_address
	wire         cpu_1f_instruction_master_read;                               // cpu_1f:i_read -> mm_interconnect_0:cpu_1f_instruction_master_read
	wire         cpu_1e_mm_bridge_0_m0_waitrequest;                            // mm_interconnect_0:CPU_1e_mm_bridge_0_m0_waitrequest -> CPU_1e:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1e_mm_bridge_0_m0_readdata;                               // mm_interconnect_0:CPU_1e_mm_bridge_0_m0_readdata -> CPU_1e:mm_bridge_0_m0_readdata
	wire         cpu_1e_mm_bridge_0_m0_debugaccess;                            // CPU_1e:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_debugaccess
	wire  [27:0] cpu_1e_mm_bridge_0_m0_address;                                // CPU_1e:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_address
	wire         cpu_1e_mm_bridge_0_m0_read;                                   // CPU_1e:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_read
	wire   [3:0] cpu_1e_mm_bridge_0_m0_byteenable;                             // CPU_1e:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_byteenable
	wire         cpu_1e_mm_bridge_0_m0_readdatavalid;                          // mm_interconnect_0:CPU_1e_mm_bridge_0_m0_readdatavalid -> CPU_1e:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1e_mm_bridge_0_m0_writedata;                              // CPU_1e:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_writedata
	wire         cpu_1e_mm_bridge_0_m0_write;                                  // CPU_1e:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_write
	wire   [0:0] cpu_1e_mm_bridge_0_m0_burstcount;                             // CPU_1e:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1e_mm_bridge_0_m0_burstcount
	wire         cpu_1d_mm_bridge_0_m0_waitrequest;                            // mm_interconnect_0:CPU_1d_mm_bridge_0_m0_waitrequest -> CPU_1d:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1d_mm_bridge_0_m0_readdata;                               // mm_interconnect_0:CPU_1d_mm_bridge_0_m0_readdata -> CPU_1d:mm_bridge_0_m0_readdata
	wire         cpu_1d_mm_bridge_0_m0_debugaccess;                            // CPU_1d:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1d_mm_bridge_0_m0_debugaccess
	wire  [27:0] cpu_1d_mm_bridge_0_m0_address;                                // CPU_1d:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1d_mm_bridge_0_m0_address
	wire         cpu_1d_mm_bridge_0_m0_read;                                   // CPU_1d:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1d_mm_bridge_0_m0_read
	wire   [3:0] cpu_1d_mm_bridge_0_m0_byteenable;                             // CPU_1d:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1d_mm_bridge_0_m0_byteenable
	wire         cpu_1d_mm_bridge_0_m0_readdatavalid;                          // mm_interconnect_0:CPU_1d_mm_bridge_0_m0_readdatavalid -> CPU_1d:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1d_mm_bridge_0_m0_writedata;                              // CPU_1d:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1d_mm_bridge_0_m0_writedata
	wire         cpu_1d_mm_bridge_0_m0_write;                                  // CPU_1d:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1d_mm_bridge_0_m0_write
	wire   [0:0] cpu_1d_mm_bridge_0_m0_burstcount;                             // CPU_1d:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1d_mm_bridge_0_m0_burstcount
	wire         cpu_1c_mm_bridge_0_m0_waitrequest;                            // mm_interconnect_0:CPU_1c_mm_bridge_0_m0_waitrequest -> CPU_1c:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1c_mm_bridge_0_m0_readdata;                               // mm_interconnect_0:CPU_1c_mm_bridge_0_m0_readdata -> CPU_1c:mm_bridge_0_m0_readdata
	wire         cpu_1c_mm_bridge_0_m0_debugaccess;                            // CPU_1c:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1c_mm_bridge_0_m0_debugaccess
	wire  [27:0] cpu_1c_mm_bridge_0_m0_address;                                // CPU_1c:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1c_mm_bridge_0_m0_address
	wire         cpu_1c_mm_bridge_0_m0_read;                                   // CPU_1c:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1c_mm_bridge_0_m0_read
	wire   [3:0] cpu_1c_mm_bridge_0_m0_byteenable;                             // CPU_1c:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1c_mm_bridge_0_m0_byteenable
	wire         cpu_1c_mm_bridge_0_m0_readdatavalid;                          // mm_interconnect_0:CPU_1c_mm_bridge_0_m0_readdatavalid -> CPU_1c:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1c_mm_bridge_0_m0_writedata;                              // CPU_1c:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1c_mm_bridge_0_m0_writedata
	wire         cpu_1c_mm_bridge_0_m0_write;                                  // CPU_1c:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1c_mm_bridge_0_m0_write
	wire   [0:0] cpu_1c_mm_bridge_0_m0_burstcount;                             // CPU_1c:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1c_mm_bridge_0_m0_burstcount
	wire         cpu_1b_mm_bridge_0_m0_waitrequest;                            // mm_interconnect_0:CPU_1b_mm_bridge_0_m0_waitrequest -> CPU_1b:mm_bridge_0_m0_waitrequest
	wire  [31:0] cpu_1b_mm_bridge_0_m0_readdata;                               // mm_interconnect_0:CPU_1b_mm_bridge_0_m0_readdata -> CPU_1b:mm_bridge_0_m0_readdata
	wire         cpu_1b_mm_bridge_0_m0_debugaccess;                            // CPU_1b:mm_bridge_0_m0_debugaccess -> mm_interconnect_0:CPU_1b_mm_bridge_0_m0_debugaccess
	wire  [27:0] cpu_1b_mm_bridge_0_m0_address;                                // CPU_1b:mm_bridge_0_m0_address -> mm_interconnect_0:CPU_1b_mm_bridge_0_m0_address
	wire         cpu_1b_mm_bridge_0_m0_read;                                   // CPU_1b:mm_bridge_0_m0_read -> mm_interconnect_0:CPU_1b_mm_bridge_0_m0_read
	wire   [3:0] cpu_1b_mm_bridge_0_m0_byteenable;                             // CPU_1b:mm_bridge_0_m0_byteenable -> mm_interconnect_0:CPU_1b_mm_bridge_0_m0_byteenable
	wire         cpu_1b_mm_bridge_0_m0_readdatavalid;                          // mm_interconnect_0:CPU_1b_mm_bridge_0_m0_readdatavalid -> CPU_1b:mm_bridge_0_m0_readdatavalid
	wire  [31:0] cpu_1b_mm_bridge_0_m0_writedata;                              // CPU_1b:mm_bridge_0_m0_writedata -> mm_interconnect_0:CPU_1b_mm_bridge_0_m0_writedata
	wire         cpu_1b_mm_bridge_0_m0_write;                                  // CPU_1b:mm_bridge_0_m0_write -> mm_interconnect_0:CPU_1b_mm_bridge_0_m0_write
	wire   [0:0] cpu_1b_mm_bridge_0_m0_burstcount;                             // CPU_1b:mm_bridge_0_m0_burstcount -> mm_interconnect_0:CPU_1b_mm_bridge_0_m0_burstcount
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;       // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;    // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sys_id_control_slave_readdata;              // sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sys_id_control_slave_address;               // mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;               // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;            // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;            // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                   // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;             // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                  // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;              // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_fifo_q_1_in_waitrequest;                    // fifo_q_1:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_1_in_waitrequest
	wire         mm_interconnect_0_fifo_q_1_in_write;                          // mm_interconnect_0:fifo_q_1_in_write -> fifo_q_1:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_1_in_writedata;                      // mm_interconnect_0:fifo_q_1_in_writedata -> fifo_q_1:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_2_in_waitrequest;                    // fifo_q_2:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_2_in_waitrequest
	wire         mm_interconnect_0_fifo_q_2_in_write;                          // mm_interconnect_0:fifo_q_2_in_write -> fifo_q_2:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_2_in_writedata;                      // mm_interconnect_0:fifo_q_2_in_writedata -> fifo_q_2:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_3_in_waitrequest;                    // fifo_q_3:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_3_in_waitrequest
	wire         mm_interconnect_0_fifo_q_3_in_write;                          // mm_interconnect_0:fifo_q_3_in_write -> fifo_q_3:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_3_in_writedata;                      // mm_interconnect_0:fifo_q_3_in_writedata -> fifo_q_3:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_4_in_waitrequest;                    // fifo_q_4:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_4_in_waitrequest
	wire         mm_interconnect_0_fifo_q_4_in_write;                          // mm_interconnect_0:fifo_q_4_in_write -> fifo_q_4:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_4_in_writedata;                      // mm_interconnect_0:fifo_q_4_in_writedata -> fifo_q_4:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_5_in_waitrequest;                    // fifo_q_5:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_5_in_waitrequest
	wire         mm_interconnect_0_fifo_q_5_in_write;                          // mm_interconnect_0:fifo_q_5_in_write -> fifo_q_5:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_5_in_writedata;                      // mm_interconnect_0:fifo_q_5_in_writedata -> fifo_q_5:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_q_6_in_waitrequest;                    // fifo_q_6:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_q_6_in_waitrequest
	wire         mm_interconnect_0_fifo_q_6_in_write;                          // mm_interconnect_0:fifo_q_6_in_write -> fifo_q_6:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_6_in_writedata;                      // mm_interconnect_0:fifo_q_6_in_writedata -> fifo_q_6:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_q_1_in_csr_readdata;                   // fifo_q_1:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_1_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_q_1_in_csr_address;                    // mm_interconnect_0:fifo_q_1_in_csr_address -> fifo_q_1:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_1_in_csr_read;                       // mm_interconnect_0:fifo_q_1_in_csr_read -> fifo_q_1:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_q_1_in_csr_write;                      // mm_interconnect_0:fifo_q_1_in_csr_write -> fifo_q_1:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_1_in_csr_writedata;                  // mm_interconnect_0:fifo_q_1_in_csr_writedata -> fifo_q_1:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_q_2_in_csr_readdata;                   // fifo_q_2:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_2_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_q_2_in_csr_address;                    // mm_interconnect_0:fifo_q_2_in_csr_address -> fifo_q_2:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_2_in_csr_read;                       // mm_interconnect_0:fifo_q_2_in_csr_read -> fifo_q_2:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_q_2_in_csr_write;                      // mm_interconnect_0:fifo_q_2_in_csr_write -> fifo_q_2:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_2_in_csr_writedata;                  // mm_interconnect_0:fifo_q_2_in_csr_writedata -> fifo_q_2:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_q_3_in_csr_readdata;                   // fifo_q_3:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_3_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_q_3_in_csr_address;                    // mm_interconnect_0:fifo_q_3_in_csr_address -> fifo_q_3:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_3_in_csr_read;                       // mm_interconnect_0:fifo_q_3_in_csr_read -> fifo_q_3:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_q_3_in_csr_write;                      // mm_interconnect_0:fifo_q_3_in_csr_write -> fifo_q_3:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_3_in_csr_writedata;                  // mm_interconnect_0:fifo_q_3_in_csr_writedata -> fifo_q_3:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_q_4_in_csr_readdata;                   // fifo_q_4:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_4_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_q_4_in_csr_address;                    // mm_interconnect_0:fifo_q_4_in_csr_address -> fifo_q_4:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_4_in_csr_read;                       // mm_interconnect_0:fifo_q_4_in_csr_read -> fifo_q_4:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_q_4_in_csr_write;                      // mm_interconnect_0:fifo_q_4_in_csr_write -> fifo_q_4:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_4_in_csr_writedata;                  // mm_interconnect_0:fifo_q_4_in_csr_writedata -> fifo_q_4:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_q_5_in_csr_readdata;                   // fifo_q_5:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_5_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_q_5_in_csr_address;                    // mm_interconnect_0:fifo_q_5_in_csr_address -> fifo_q_5:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_5_in_csr_read;                       // mm_interconnect_0:fifo_q_5_in_csr_read -> fifo_q_5:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_q_5_in_csr_write;                      // mm_interconnect_0:fifo_q_5_in_csr_write -> fifo_q_5:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_5_in_csr_writedata;                  // mm_interconnect_0:fifo_q_5_in_csr_writedata -> fifo_q_5:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_q_6_in_csr_readdata;                   // fifo_q_6:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_q_6_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_q_6_in_csr_address;                    // mm_interconnect_0:fifo_q_6_in_csr_address -> fifo_q_6:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_q_6_in_csr_read;                       // mm_interconnect_0:fifo_q_6_in_csr_read -> fifo_q_6:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_q_6_in_csr_write;                      // mm_interconnect_0:fifo_q_6_in_csr_write -> fifo_q_6:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_q_6_in_csr_writedata;                  // mm_interconnect_0:fifo_q_6_in_csr_writedata -> fifo_q_6:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                     // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                      // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                         // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                        // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                    // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;             // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;               // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;            // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;                // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;                   // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;             // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;          // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;                  // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;              // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         mm_interconnect_0_timer_s1_chipselect;                        // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                          // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                           // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                             // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                         // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire  [31:0] mm_interconnect_0_cpu_1f_debug_mem_slave_readdata;            // cpu_1f:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1f_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_1f_debug_mem_slave_waitrequest;         // cpu_1f:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1f_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_1f_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_1f_debug_mem_slave_debugaccess -> cpu_1f:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_1f_debug_mem_slave_address;             // mm_interconnect_0:cpu_1f_debug_mem_slave_address -> cpu_1f:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_1f_debug_mem_slave_read;                // mm_interconnect_0:cpu_1f_debug_mem_slave_read -> cpu_1f:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_1f_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_1f_debug_mem_slave_byteenable -> cpu_1f:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_1f_debug_mem_slave_write;               // mm_interconnect_0:cpu_1f_debug_mem_slave_write -> cpu_1f:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_1f_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_1f_debug_mem_slave_writedata -> cpu_1f:debug_mem_slave_writedata
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_chipselect -> jtag_uart_1f:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_readdata;    // jtag_uart_1f:av_readdata -> mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_waitrequest; // jtag_uart_1f:av_waitrequest -> mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_address -> jtag_uart_1f:av_address
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_read -> jtag_uart_1f:av_read_n
	wire         mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_write -> jtag_uart_1f:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1f_avalon_jtag_slave_writedata -> jtag_uart_1f:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_1f_control_slave_readdata;            // sysid_1f:readdata -> mm_interconnect_0:sysid_1f_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_1f_control_slave_address;             // mm_interconnect_0:sysid_1f_control_slave_address -> sysid_1f:address
	wire  [31:0] mm_interconnect_0_fifo_1e_in_csr_readdata;                    // fifo_1e:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_1e_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_1e_in_csr_address;                     // mm_interconnect_0:fifo_1e_in_csr_address -> fifo_1e:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_1e_in_csr_read;                        // mm_interconnect_0:fifo_1e_in_csr_read -> fifo_1e:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_1e_in_csr_write;                       // mm_interconnect_0:fifo_1e_in_csr_write -> fifo_1e:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_1e_in_csr_writedata;                   // mm_interconnect_0:fifo_1e_in_csr_writedata -> fifo_1e:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_1e_out_readdata;                       // fifo_1e:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_1e_out_readdata
	wire         mm_interconnect_0_fifo_1e_out_waitrequest;                    // fifo_1e:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_1e_out_waitrequest
	wire         mm_interconnect_0_fifo_1e_out_read;                           // mm_interconnect_0:fifo_1e_out_read -> fifo_1e:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_6_out_readdata;                      // fifo_q_6:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_6_out_readdata
	wire         mm_interconnect_0_fifo_q_6_out_waitrequest;                   // fifo_q_6:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_6_out_waitrequest
	wire         mm_interconnect_0_fifo_q_6_out_read;                          // mm_interconnect_0:fifo_q_6_out_read -> fifo_q_6:avalonmm_read_slave_read
	wire         mm_interconnect_0_timer_1f_s1_chipselect;                     // mm_interconnect_0:timer_1f_s1_chipselect -> timer_1f:chipselect
	wire  [15:0] mm_interconnect_0_timer_1f_s1_readdata;                       // timer_1f:readdata -> mm_interconnect_0:timer_1f_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1f_s1_address;                        // mm_interconnect_0:timer_1f_s1_address -> timer_1f:address
	wire         mm_interconnect_0_timer_1f_s1_write;                          // mm_interconnect_0:timer_1f_s1_write -> timer_1f:write_n
	wire  [15:0] mm_interconnect_0_timer_1f_s1_writedata;                      // mm_interconnect_0:timer_1f_s1_writedata -> timer_1f:writedata
	wire         mm_interconnect_0_fifo_1e_in_waitrequest;                     // fifo_1e:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_1e_in_waitrequest
	wire         mm_interconnect_0_fifo_1e_in_write;                           // mm_interconnect_0:fifo_1e_in_write -> fifo_1e:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_1e_in_writedata;                       // mm_interconnect_0:fifo_1e_in_writedata -> fifo_1e:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_1d_in_csr_readdata;                    // fifo_1d:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_1d_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_1d_in_csr_address;                     // mm_interconnect_0:fifo_1d_in_csr_address -> fifo_1d:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_1d_in_csr_read;                        // mm_interconnect_0:fifo_1d_in_csr_read -> fifo_1d:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_1d_in_csr_write;                       // mm_interconnect_0:fifo_1d_in_csr_write -> fifo_1d:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_1d_in_csr_writedata;                   // mm_interconnect_0:fifo_1d_in_csr_writedata -> fifo_1d:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_1d_out_readdata;                       // fifo_1d:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_1d_out_readdata
	wire         mm_interconnect_0_fifo_1d_out_waitrequest;                    // fifo_1d:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_1d_out_waitrequest
	wire         mm_interconnect_0_fifo_1d_out_read;                           // mm_interconnect_0:fifo_1d_out_read -> fifo_1d:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_5_out_readdata;                      // fifo_q_5:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_5_out_readdata
	wire         mm_interconnect_0_fifo_q_5_out_waitrequest;                   // fifo_q_5:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_5_out_waitrequest
	wire         mm_interconnect_0_fifo_q_5_out_read;                          // mm_interconnect_0:fifo_q_5_out_read -> fifo_q_5:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_1d_in_waitrequest;                     // fifo_1d:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_1d_in_waitrequest
	wire         mm_interconnect_0_fifo_1d_in_write;                           // mm_interconnect_0:fifo_1d_in_write -> fifo_1d:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_1d_in_writedata;                       // mm_interconnect_0:fifo_1d_in_writedata -> fifo_1d:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_1c_in_csr_readdata;                    // fifo_1c:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_1c_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_1c_in_csr_address;                     // mm_interconnect_0:fifo_1c_in_csr_address -> fifo_1c:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_1c_in_csr_read;                        // mm_interconnect_0:fifo_1c_in_csr_read -> fifo_1c:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_1c_in_csr_write;                       // mm_interconnect_0:fifo_1c_in_csr_write -> fifo_1c:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_1c_in_csr_writedata;                   // mm_interconnect_0:fifo_1c_in_csr_writedata -> fifo_1c:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_1c_out_readdata;                       // fifo_1c:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_1c_out_readdata
	wire         mm_interconnect_0_fifo_1c_out_waitrequest;                    // fifo_1c:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_1c_out_waitrequest
	wire         mm_interconnect_0_fifo_1c_out_read;                           // mm_interconnect_0:fifo_1c_out_read -> fifo_1c:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_4_out_readdata;                      // fifo_q_4:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_4_out_readdata
	wire         mm_interconnect_0_fifo_q_4_out_waitrequest;                   // fifo_q_4:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_4_out_waitrequest
	wire         mm_interconnect_0_fifo_q_4_out_read;                          // mm_interconnect_0:fifo_q_4_out_read -> fifo_q_4:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_1c_in_waitrequest;                     // fifo_1c:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_1c_in_waitrequest
	wire         mm_interconnect_0_fifo_1c_in_write;                           // mm_interconnect_0:fifo_1c_in_write -> fifo_1c:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_1c_in_writedata;                       // mm_interconnect_0:fifo_1c_in_writedata -> fifo_1c:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_1b_in_csr_readdata;                    // fifo_1b:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_1b_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_1b_in_csr_address;                     // mm_interconnect_0:fifo_1b_in_csr_address -> fifo_1b:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_1b_in_csr_read;                        // mm_interconnect_0:fifo_1b_in_csr_read -> fifo_1b:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_1b_in_csr_write;                       // mm_interconnect_0:fifo_1b_in_csr_write -> fifo_1b:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_1b_in_csr_writedata;                   // mm_interconnect_0:fifo_1b_in_csr_writedata -> fifo_1b:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_1b_out_readdata;                       // fifo_1b:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_1b_out_readdata
	wire         mm_interconnect_0_fifo_1b_out_waitrequest;                    // fifo_1b:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_1b_out_waitrequest
	wire         mm_interconnect_0_fifo_1b_out_read;                           // mm_interconnect_0:fifo_1b_out_read -> fifo_1b:avalonmm_read_slave_read
	wire         mm_interconnect_0_fifo_1b_in_waitrequest;                     // fifo_1b:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_1b_in_waitrequest
	wire         mm_interconnect_0_fifo_1b_in_write;                           // mm_interconnect_0:fifo_1b_in_write -> fifo_1b:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_1b_in_writedata;                       // mm_interconnect_0:fifo_1b_in_writedata -> fifo_1b:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_fifo_q_1_out_readdata;                      // fifo_q_1:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_1_out_readdata
	wire         mm_interconnect_0_fifo_q_1_out_waitrequest;                   // fifo_q_1:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_1_out_waitrequest
	wire         mm_interconnect_0_fifo_q_1_out_read;                          // mm_interconnect_0:fifo_q_1_out_read -> fifo_q_1:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_2_out_readdata;                      // fifo_q_2:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_2_out_readdata
	wire         mm_interconnect_0_fifo_q_2_out_waitrequest;                   // fifo_q_2:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_2_out_waitrequest
	wire         mm_interconnect_0_fifo_q_2_out_read;                          // mm_interconnect_0:fifo_q_2_out_read -> fifo_q_2:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_q_3_out_readdata;                      // fifo_q_3:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_q_3_out_readdata
	wire         mm_interconnect_0_fifo_q_3_out_waitrequest;                   // fifo_q_3:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_q_3_out_waitrequest
	wire         mm_interconnect_0_fifo_q_3_out_read;                          // mm_interconnect_0:fifo_q_3_out_read -> fifo_q_3:avalonmm_read_slave_read
	wire         irq_mapper_receiver0_irq;                                     // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                                  // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_001_receiver0_irq;                                 // timer_1f:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                 // jtag_uart_1f:av_irq -> irq_mapper_001:receiver1_irq
	wire  [31:0] cpu_1f_irq_irq;                                               // irq_mapper_001:sender_irq -> cpu_1f:irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [CPU_1b:reset_bridge_0_in_reset_reset, CPU_1c:reset_bridge_0_in_reset_reset, CPU_1d:reset_bridge_0_in_reset_reset, CPU_1e:reset_bridge_0_in_reset_reset, mm_interconnect_0:CPU_1e_reset_bridge_0_in_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [cpu:reset_n, cpu_1f:reset_n, fifo_1b:reset_n, fifo_1c:reset_n, fifo_1d:reset_n, fifo_1e:reset_n, fifo_q_1:reset_n, fifo_q_2:reset_n, fifo_q_3:reset_n, fifo_q_4:reset_n, fifo_q_5:reset_n, fifo_q_6:reset_n, irq_mapper:reset, irq_mapper_001:reset, jtag_uart:rst_n, jtag_uart_1f:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram_controller:reset_n, sys_id:reset_n, sysid_1f:reset_n, timer:reset_n, timer_1f:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                       // rst_controller_001:reset_req -> [cpu:reset_req, cpu_1f:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                // cpu:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         cpu_1f_debug_reset_request_reset;                             // cpu_1f:debug_reset_request -> [rst_controller_001:reset_in2, rst_controller_002:reset_in2]
	wire         rst_controller_002_reset_out_reset;                           // rst_controller_002:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	TOP_MSOC_CPU_1b cpu_1b (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                          //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1b_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1b_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1b_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1b_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1b_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1b_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1b_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1b_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1b_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1b_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)       // reset_bridge_0_in_reset.reset
	);

	TOP_MSOC_CPU_1c cpu_1c (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                          //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1c_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1c_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1c_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1c_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1c_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1c_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1c_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1c_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1c_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1c_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)       // reset_bridge_0_in_reset.reset
	);

	TOP_MSOC_CPU_1d cpu_1d (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                          //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1d_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1d_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1d_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1d_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1d_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1d_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1d_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1d_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1d_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1d_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)       // reset_bridge_0_in_reset.reset
	);

	TOP_MSOC_CPU_1e cpu_1e (
		.clock_bridge_0_in_clk_clk     (pll_c0_clk),                          //   clock_bridge_0_in_clk.clk
		.mm_bridge_0_m0_waitrequest    (cpu_1e_mm_bridge_0_m0_waitrequest),   //          mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata       (cpu_1e_mm_bridge_0_m0_readdata),      //                        .readdata
		.mm_bridge_0_m0_readdatavalid  (cpu_1e_mm_bridge_0_m0_readdatavalid), //                        .readdatavalid
		.mm_bridge_0_m0_burstcount     (cpu_1e_mm_bridge_0_m0_burstcount),    //                        .burstcount
		.mm_bridge_0_m0_writedata      (cpu_1e_mm_bridge_0_m0_writedata),     //                        .writedata
		.mm_bridge_0_m0_address        (cpu_1e_mm_bridge_0_m0_address),       //                        .address
		.mm_bridge_0_m0_write          (cpu_1e_mm_bridge_0_m0_write),         //                        .write
		.mm_bridge_0_m0_read           (cpu_1e_mm_bridge_0_m0_read),          //                        .read
		.mm_bridge_0_m0_byteenable     (cpu_1e_mm_bridge_0_m0_byteenable),    //                        .byteenable
		.mm_bridge_0_m0_debugaccess    (cpu_1e_mm_bridge_0_m0_debugaccess),   //                        .debugaccess
		.reset_bridge_0_in_reset_reset (rst_controller_reset_out_reset)       // reset_bridge_0_in_reset.reset
	);

	TOP_MSOC_cpu cpu (
		.clk                                 (pll_c0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	TOP_MSOC_cpu_1f cpu_1f (
		.clk                                 (pll_c0_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                  //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),               //                          .reset_req
		.d_address                           (cpu_1f_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_1f_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_1f_data_master_read),                              //                          .read
		.d_readdata                          (cpu_1f_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_1f_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_1f_data_master_write),                             //                          .write
		.d_writedata                         (cpu_1f_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_1f_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_1f_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_1f_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_1f_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_1f_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_1f_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_1f_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_1f_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_1f_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_1f_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_1f_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_1f_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_1f_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_1f_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_1f_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	TOP_MSOC_fifo_1b fifo_1b (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_1b_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_1b_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_1b_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_1b_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_1b_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_1b_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_1b_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_1b_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_1b_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_1b_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_1b_in_csr_readdata)   //         .readdata
	);

	TOP_MSOC_fifo_1b fifo_1c (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_1c_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_1c_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_1c_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_1c_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_1c_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_1c_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_1c_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_1c_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_1c_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_1c_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_1c_in_csr_readdata)   //         .readdata
	);

	TOP_MSOC_fifo_1b fifo_1d (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_1d_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_1d_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_1d_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_1d_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_1d_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_1d_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_1d_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_1d_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_1d_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_1d_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_1d_in_csr_readdata)   //         .readdata
	);

	TOP_MSOC_fifo_1b fifo_1e (
		.wrclock                          (pll_c0_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),        // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_1e_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_1e_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_1e_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_1e_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_1e_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_1e_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_1e_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_1e_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_1e_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_1e_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_1e_in_csr_readdata)   //         .readdata
	);

	TOP_MSOC_fifo_q_1 fifo_q_1 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_1_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_1_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_1_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_1_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_1_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_1_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_1_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_1_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_1_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_1_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_1_in_csr_readdata)   //         .readdata
	);

	TOP_MSOC_fifo_q_1 fifo_q_2 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_2_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_2_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_2_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_2_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_2_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_2_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_2_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_2_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_2_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_2_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_2_in_csr_readdata)   //         .readdata
	);

	TOP_MSOC_fifo_q_1 fifo_q_3 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_3_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_3_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_3_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_3_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_3_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_3_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_3_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_3_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_3_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_3_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_3_in_csr_readdata)   //         .readdata
	);

	TOP_MSOC_fifo_1b fifo_q_4 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_4_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_4_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_4_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_4_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_4_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_4_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_4_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_4_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_4_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_4_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_4_in_csr_readdata)   //         .readdata
	);

	TOP_MSOC_fifo_1b fifo_q_5 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_5_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_5_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_5_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_5_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_5_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_5_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_5_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_5_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_5_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_5_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_5_in_csr_readdata)   //         .readdata
	);

	TOP_MSOC_fifo_1b fifo_q_6 (
		.wrclock                          (pll_c0_clk),                                  //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_q_6_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_q_6_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_q_6_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_q_6_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_q_6_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_q_6_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_q_6_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_q_6_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_q_6_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_q_6_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_q_6_in_csr_readdata)   //         .readdata
	);

	TOP_MSOC_jtag_uart jtag_uart (
		.clk            (pll_c0_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	TOP_MSOC_jtag_uart jtag_uart_1f (
		.clk            (pll_c0_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                          //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver1_irq)                                  //               irq.irq
	);

	TOP_MSOC_pll pll (
		.clk                (clk_clk),                                   //       inclk_interface.clk
		.reset              (rst_controller_002_reset_out_reset),        // inclk_interface_reset.reset
		.read               (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0                 (pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                             //                    c1.clk
		.scandone           (),                                          //           (terminated)
		.scandataout        (),                                          //           (terminated)
		.phasecounterselect (4'b0000),                                   //           (terminated)
		.phaseupdown        (1'b0),                                      //           (terminated)
		.phasestep          (1'b0),                                      //           (terminated)
		.scanclk            (1'b0),                                      //           (terminated)
		.scanclkena         (1'b0),                                      //           (terminated)
		.scandata           (1'b0),                                      //           (terminated)
		.configupdate       (1'b0),                                      //           (terminated)
		.areset             (1'b0),                                      //           (terminated)
		.locked             (),                                          //           (terminated)
		.phasedone          ()                                           //           (terminated)
	);

	TOP_MSOC_sdram_controller sdram_controller (
		.clk            (pll_c0_clk),                                          //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                 // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                           //      .export
	);

	TOP_MSOC_sys_id sys_id (
		.clock    (pll_c0_clk),                                      //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),             //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //              .address
	);

	TOP_MSOC_sysid_1f sysid_1f (
		.clock    (pll_c0_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),               //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_1f_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_1f_control_slave_address)   //              .address
	);

	TOP_MSOC_timer timer (
		.clk        (pll_c0_clk),                            //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	TOP_MSOC_timer timer_1f (
		.clk        (pll_c0_clk),                               //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.address    (mm_interconnect_0_timer_1f_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1f_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1f_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1f_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1f_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver0_irq)              //   irq.irq
	);

	TOP_MSOC_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                              (clk_clk),                                                      //                                            clock_clk.clk
		.pll_c0_clk                                                 (pll_c0_clk),                                                   //                                               pll_c0.clk
		.CPU_1e_reset_bridge_0_in_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // CPU_1e_reset_bridge_0_in_reset_reset_bridge_in_reset.reset
		.cpu_reset_reset_bridge_in_reset_reset                      (rst_controller_001_reset_out_reset),                           //                      cpu_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset      (rst_controller_002_reset_out_reset),                           //      pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                    (cpu_data_master_address),                                      //                                      cpu_data_master.address
		.cpu_data_master_waitrequest                                (cpu_data_master_waitrequest),                                  //                                                     .waitrequest
		.cpu_data_master_byteenable                                 (cpu_data_master_byteenable),                                   //                                                     .byteenable
		.cpu_data_master_read                                       (cpu_data_master_read),                                         //                                                     .read
		.cpu_data_master_readdata                                   (cpu_data_master_readdata),                                     //                                                     .readdata
		.cpu_data_master_write                                      (cpu_data_master_write),                                        //                                                     .write
		.cpu_data_master_writedata                                  (cpu_data_master_writedata),                                    //                                                     .writedata
		.cpu_data_master_debugaccess                                (cpu_data_master_debugaccess),                                  //                                                     .debugaccess
		.cpu_instruction_master_address                             (cpu_instruction_master_address),                               //                               cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                         (cpu_instruction_master_waitrequest),                           //                                                     .waitrequest
		.cpu_instruction_master_read                                (cpu_instruction_master_read),                                  //                                                     .read
		.cpu_instruction_master_readdata                            (cpu_instruction_master_readdata),                              //                                                     .readdata
		.CPU_1b_mm_bridge_0_m0_address                              (cpu_1b_mm_bridge_0_m0_address),                                //                                CPU_1b_mm_bridge_0_m0.address
		.CPU_1b_mm_bridge_0_m0_waitrequest                          (cpu_1b_mm_bridge_0_m0_waitrequest),                            //                                                     .waitrequest
		.CPU_1b_mm_bridge_0_m0_burstcount                           (cpu_1b_mm_bridge_0_m0_burstcount),                             //                                                     .burstcount
		.CPU_1b_mm_bridge_0_m0_byteenable                           (cpu_1b_mm_bridge_0_m0_byteenable),                             //                                                     .byteenable
		.CPU_1b_mm_bridge_0_m0_read                                 (cpu_1b_mm_bridge_0_m0_read),                                   //                                                     .read
		.CPU_1b_mm_bridge_0_m0_readdata                             (cpu_1b_mm_bridge_0_m0_readdata),                               //                                                     .readdata
		.CPU_1b_mm_bridge_0_m0_readdatavalid                        (cpu_1b_mm_bridge_0_m0_readdatavalid),                          //                                                     .readdatavalid
		.CPU_1b_mm_bridge_0_m0_write                                (cpu_1b_mm_bridge_0_m0_write),                                  //                                                     .write
		.CPU_1b_mm_bridge_0_m0_writedata                            (cpu_1b_mm_bridge_0_m0_writedata),                              //                                                     .writedata
		.CPU_1b_mm_bridge_0_m0_debugaccess                          (cpu_1b_mm_bridge_0_m0_debugaccess),                            //                                                     .debugaccess
		.CPU_1c_mm_bridge_0_m0_address                              (cpu_1c_mm_bridge_0_m0_address),                                //                                CPU_1c_mm_bridge_0_m0.address
		.CPU_1c_mm_bridge_0_m0_waitrequest                          (cpu_1c_mm_bridge_0_m0_waitrequest),                            //                                                     .waitrequest
		.CPU_1c_mm_bridge_0_m0_burstcount                           (cpu_1c_mm_bridge_0_m0_burstcount),                             //                                                     .burstcount
		.CPU_1c_mm_bridge_0_m0_byteenable                           (cpu_1c_mm_bridge_0_m0_byteenable),                             //                                                     .byteenable
		.CPU_1c_mm_bridge_0_m0_read                                 (cpu_1c_mm_bridge_0_m0_read),                                   //                                                     .read
		.CPU_1c_mm_bridge_0_m0_readdata                             (cpu_1c_mm_bridge_0_m0_readdata),                               //                                                     .readdata
		.CPU_1c_mm_bridge_0_m0_readdatavalid                        (cpu_1c_mm_bridge_0_m0_readdatavalid),                          //                                                     .readdatavalid
		.CPU_1c_mm_bridge_0_m0_write                                (cpu_1c_mm_bridge_0_m0_write),                                  //                                                     .write
		.CPU_1c_mm_bridge_0_m0_writedata                            (cpu_1c_mm_bridge_0_m0_writedata),                              //                                                     .writedata
		.CPU_1c_mm_bridge_0_m0_debugaccess                          (cpu_1c_mm_bridge_0_m0_debugaccess),                            //                                                     .debugaccess
		.CPU_1d_mm_bridge_0_m0_address                              (cpu_1d_mm_bridge_0_m0_address),                                //                                CPU_1d_mm_bridge_0_m0.address
		.CPU_1d_mm_bridge_0_m0_waitrequest                          (cpu_1d_mm_bridge_0_m0_waitrequest),                            //                                                     .waitrequest
		.CPU_1d_mm_bridge_0_m0_burstcount                           (cpu_1d_mm_bridge_0_m0_burstcount),                             //                                                     .burstcount
		.CPU_1d_mm_bridge_0_m0_byteenable                           (cpu_1d_mm_bridge_0_m0_byteenable),                             //                                                     .byteenable
		.CPU_1d_mm_bridge_0_m0_read                                 (cpu_1d_mm_bridge_0_m0_read),                                   //                                                     .read
		.CPU_1d_mm_bridge_0_m0_readdata                             (cpu_1d_mm_bridge_0_m0_readdata),                               //                                                     .readdata
		.CPU_1d_mm_bridge_0_m0_readdatavalid                        (cpu_1d_mm_bridge_0_m0_readdatavalid),                          //                                                     .readdatavalid
		.CPU_1d_mm_bridge_0_m0_write                                (cpu_1d_mm_bridge_0_m0_write),                                  //                                                     .write
		.CPU_1d_mm_bridge_0_m0_writedata                            (cpu_1d_mm_bridge_0_m0_writedata),                              //                                                     .writedata
		.CPU_1d_mm_bridge_0_m0_debugaccess                          (cpu_1d_mm_bridge_0_m0_debugaccess),                            //                                                     .debugaccess
		.CPU_1e_mm_bridge_0_m0_address                              (cpu_1e_mm_bridge_0_m0_address),                                //                                CPU_1e_mm_bridge_0_m0.address
		.CPU_1e_mm_bridge_0_m0_waitrequest                          (cpu_1e_mm_bridge_0_m0_waitrequest),                            //                                                     .waitrequest
		.CPU_1e_mm_bridge_0_m0_burstcount                           (cpu_1e_mm_bridge_0_m0_burstcount),                             //                                                     .burstcount
		.CPU_1e_mm_bridge_0_m0_byteenable                           (cpu_1e_mm_bridge_0_m0_byteenable),                             //                                                     .byteenable
		.CPU_1e_mm_bridge_0_m0_read                                 (cpu_1e_mm_bridge_0_m0_read),                                   //                                                     .read
		.CPU_1e_mm_bridge_0_m0_readdata                             (cpu_1e_mm_bridge_0_m0_readdata),                               //                                                     .readdata
		.CPU_1e_mm_bridge_0_m0_readdatavalid                        (cpu_1e_mm_bridge_0_m0_readdatavalid),                          //                                                     .readdatavalid
		.CPU_1e_mm_bridge_0_m0_write                                (cpu_1e_mm_bridge_0_m0_write),                                  //                                                     .write
		.CPU_1e_mm_bridge_0_m0_writedata                            (cpu_1e_mm_bridge_0_m0_writedata),                              //                                                     .writedata
		.CPU_1e_mm_bridge_0_m0_debugaccess                          (cpu_1e_mm_bridge_0_m0_debugaccess),                            //                                                     .debugaccess
		.cpu_1f_data_master_address                                 (cpu_1f_data_master_address),                                   //                                   cpu_1f_data_master.address
		.cpu_1f_data_master_waitrequest                             (cpu_1f_data_master_waitrequest),                               //                                                     .waitrequest
		.cpu_1f_data_master_byteenable                              (cpu_1f_data_master_byteenable),                                //                                                     .byteenable
		.cpu_1f_data_master_read                                    (cpu_1f_data_master_read),                                      //                                                     .read
		.cpu_1f_data_master_readdata                                (cpu_1f_data_master_readdata),                                  //                                                     .readdata
		.cpu_1f_data_master_write                                   (cpu_1f_data_master_write),                                     //                                                     .write
		.cpu_1f_data_master_writedata                               (cpu_1f_data_master_writedata),                                 //                                                     .writedata
		.cpu_1f_data_master_debugaccess                             (cpu_1f_data_master_debugaccess),                               //                                                     .debugaccess
		.cpu_1f_instruction_master_address                          (cpu_1f_instruction_master_address),                            //                            cpu_1f_instruction_master.address
		.cpu_1f_instruction_master_waitrequest                      (cpu_1f_instruction_master_waitrequest),                        //                                                     .waitrequest
		.cpu_1f_instruction_master_read                             (cpu_1f_instruction_master_read),                               //                                                     .read
		.cpu_1f_instruction_master_readdata                         (cpu_1f_instruction_master_readdata),                           //                                                     .readdata
		.cpu_debug_mem_slave_address                                (mm_interconnect_0_cpu_debug_mem_slave_address),                //                                  cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                  (mm_interconnect_0_cpu_debug_mem_slave_write),                  //                                                     .write
		.cpu_debug_mem_slave_read                                   (mm_interconnect_0_cpu_debug_mem_slave_read),                   //                                                     .read
		.cpu_debug_mem_slave_readdata                               (mm_interconnect_0_cpu_debug_mem_slave_readdata),               //                                                     .readdata
		.cpu_debug_mem_slave_writedata                              (mm_interconnect_0_cpu_debug_mem_slave_writedata),              //                                                     .writedata
		.cpu_debug_mem_slave_byteenable                             (mm_interconnect_0_cpu_debug_mem_slave_byteenable),             //                                                     .byteenable
		.cpu_debug_mem_slave_waitrequest                            (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),            //                                                     .waitrequest
		.cpu_debug_mem_slave_debugaccess                            (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),            //                                                     .debugaccess
		.cpu_1f_debug_mem_slave_address                             (mm_interconnect_0_cpu_1f_debug_mem_slave_address),             //                               cpu_1f_debug_mem_slave.address
		.cpu_1f_debug_mem_slave_write                               (mm_interconnect_0_cpu_1f_debug_mem_slave_write),               //                                                     .write
		.cpu_1f_debug_mem_slave_read                                (mm_interconnect_0_cpu_1f_debug_mem_slave_read),                //                                                     .read
		.cpu_1f_debug_mem_slave_readdata                            (mm_interconnect_0_cpu_1f_debug_mem_slave_readdata),            //                                                     .readdata
		.cpu_1f_debug_mem_slave_writedata                           (mm_interconnect_0_cpu_1f_debug_mem_slave_writedata),           //                                                     .writedata
		.cpu_1f_debug_mem_slave_byteenable                          (mm_interconnect_0_cpu_1f_debug_mem_slave_byteenable),          //                                                     .byteenable
		.cpu_1f_debug_mem_slave_waitrequest                         (mm_interconnect_0_cpu_1f_debug_mem_slave_waitrequest),         //                                                     .waitrequest
		.cpu_1f_debug_mem_slave_debugaccess                         (mm_interconnect_0_cpu_1f_debug_mem_slave_debugaccess),         //                                                     .debugaccess
		.fifo_1b_in_write                                           (mm_interconnect_0_fifo_1b_in_write),                           //                                           fifo_1b_in.write
		.fifo_1b_in_writedata                                       (mm_interconnect_0_fifo_1b_in_writedata),                       //                                                     .writedata
		.fifo_1b_in_waitrequest                                     (mm_interconnect_0_fifo_1b_in_waitrequest),                     //                                                     .waitrequest
		.fifo_1b_in_csr_address                                     (mm_interconnect_0_fifo_1b_in_csr_address),                     //                                       fifo_1b_in_csr.address
		.fifo_1b_in_csr_write                                       (mm_interconnect_0_fifo_1b_in_csr_write),                       //                                                     .write
		.fifo_1b_in_csr_read                                        (mm_interconnect_0_fifo_1b_in_csr_read),                        //                                                     .read
		.fifo_1b_in_csr_readdata                                    (mm_interconnect_0_fifo_1b_in_csr_readdata),                    //                                                     .readdata
		.fifo_1b_in_csr_writedata                                   (mm_interconnect_0_fifo_1b_in_csr_writedata),                   //                                                     .writedata
		.fifo_1b_out_read                                           (mm_interconnect_0_fifo_1b_out_read),                           //                                          fifo_1b_out.read
		.fifo_1b_out_readdata                                       (mm_interconnect_0_fifo_1b_out_readdata),                       //                                                     .readdata
		.fifo_1b_out_waitrequest                                    (mm_interconnect_0_fifo_1b_out_waitrequest),                    //                                                     .waitrequest
		.fifo_1c_in_write                                           (mm_interconnect_0_fifo_1c_in_write),                           //                                           fifo_1c_in.write
		.fifo_1c_in_writedata                                       (mm_interconnect_0_fifo_1c_in_writedata),                       //                                                     .writedata
		.fifo_1c_in_waitrequest                                     (mm_interconnect_0_fifo_1c_in_waitrequest),                     //                                                     .waitrequest
		.fifo_1c_in_csr_address                                     (mm_interconnect_0_fifo_1c_in_csr_address),                     //                                       fifo_1c_in_csr.address
		.fifo_1c_in_csr_write                                       (mm_interconnect_0_fifo_1c_in_csr_write),                       //                                                     .write
		.fifo_1c_in_csr_read                                        (mm_interconnect_0_fifo_1c_in_csr_read),                        //                                                     .read
		.fifo_1c_in_csr_readdata                                    (mm_interconnect_0_fifo_1c_in_csr_readdata),                    //                                                     .readdata
		.fifo_1c_in_csr_writedata                                   (mm_interconnect_0_fifo_1c_in_csr_writedata),                   //                                                     .writedata
		.fifo_1c_out_read                                           (mm_interconnect_0_fifo_1c_out_read),                           //                                          fifo_1c_out.read
		.fifo_1c_out_readdata                                       (mm_interconnect_0_fifo_1c_out_readdata),                       //                                                     .readdata
		.fifo_1c_out_waitrequest                                    (mm_interconnect_0_fifo_1c_out_waitrequest),                    //                                                     .waitrequest
		.fifo_1d_in_write                                           (mm_interconnect_0_fifo_1d_in_write),                           //                                           fifo_1d_in.write
		.fifo_1d_in_writedata                                       (mm_interconnect_0_fifo_1d_in_writedata),                       //                                                     .writedata
		.fifo_1d_in_waitrequest                                     (mm_interconnect_0_fifo_1d_in_waitrequest),                     //                                                     .waitrequest
		.fifo_1d_in_csr_address                                     (mm_interconnect_0_fifo_1d_in_csr_address),                     //                                       fifo_1d_in_csr.address
		.fifo_1d_in_csr_write                                       (mm_interconnect_0_fifo_1d_in_csr_write),                       //                                                     .write
		.fifo_1d_in_csr_read                                        (mm_interconnect_0_fifo_1d_in_csr_read),                        //                                                     .read
		.fifo_1d_in_csr_readdata                                    (mm_interconnect_0_fifo_1d_in_csr_readdata),                    //                                                     .readdata
		.fifo_1d_in_csr_writedata                                   (mm_interconnect_0_fifo_1d_in_csr_writedata),                   //                                                     .writedata
		.fifo_1d_out_read                                           (mm_interconnect_0_fifo_1d_out_read),                           //                                          fifo_1d_out.read
		.fifo_1d_out_readdata                                       (mm_interconnect_0_fifo_1d_out_readdata),                       //                                                     .readdata
		.fifo_1d_out_waitrequest                                    (mm_interconnect_0_fifo_1d_out_waitrequest),                    //                                                     .waitrequest
		.fifo_1e_in_write                                           (mm_interconnect_0_fifo_1e_in_write),                           //                                           fifo_1e_in.write
		.fifo_1e_in_writedata                                       (mm_interconnect_0_fifo_1e_in_writedata),                       //                                                     .writedata
		.fifo_1e_in_waitrequest                                     (mm_interconnect_0_fifo_1e_in_waitrequest),                     //                                                     .waitrequest
		.fifo_1e_in_csr_address                                     (mm_interconnect_0_fifo_1e_in_csr_address),                     //                                       fifo_1e_in_csr.address
		.fifo_1e_in_csr_write                                       (mm_interconnect_0_fifo_1e_in_csr_write),                       //                                                     .write
		.fifo_1e_in_csr_read                                        (mm_interconnect_0_fifo_1e_in_csr_read),                        //                                                     .read
		.fifo_1e_in_csr_readdata                                    (mm_interconnect_0_fifo_1e_in_csr_readdata),                    //                                                     .readdata
		.fifo_1e_in_csr_writedata                                   (mm_interconnect_0_fifo_1e_in_csr_writedata),                   //                                                     .writedata
		.fifo_1e_out_read                                           (mm_interconnect_0_fifo_1e_out_read),                           //                                          fifo_1e_out.read
		.fifo_1e_out_readdata                                       (mm_interconnect_0_fifo_1e_out_readdata),                       //                                                     .readdata
		.fifo_1e_out_waitrequest                                    (mm_interconnect_0_fifo_1e_out_waitrequest),                    //                                                     .waitrequest
		.fifo_q_1_in_write                                          (mm_interconnect_0_fifo_q_1_in_write),                          //                                          fifo_q_1_in.write
		.fifo_q_1_in_writedata                                      (mm_interconnect_0_fifo_q_1_in_writedata),                      //                                                     .writedata
		.fifo_q_1_in_waitrequest                                    (mm_interconnect_0_fifo_q_1_in_waitrequest),                    //                                                     .waitrequest
		.fifo_q_1_in_csr_address                                    (mm_interconnect_0_fifo_q_1_in_csr_address),                    //                                      fifo_q_1_in_csr.address
		.fifo_q_1_in_csr_write                                      (mm_interconnect_0_fifo_q_1_in_csr_write),                      //                                                     .write
		.fifo_q_1_in_csr_read                                       (mm_interconnect_0_fifo_q_1_in_csr_read),                       //                                                     .read
		.fifo_q_1_in_csr_readdata                                   (mm_interconnect_0_fifo_q_1_in_csr_readdata),                   //                                                     .readdata
		.fifo_q_1_in_csr_writedata                                  (mm_interconnect_0_fifo_q_1_in_csr_writedata),                  //                                                     .writedata
		.fifo_q_1_out_read                                          (mm_interconnect_0_fifo_q_1_out_read),                          //                                         fifo_q_1_out.read
		.fifo_q_1_out_readdata                                      (mm_interconnect_0_fifo_q_1_out_readdata),                      //                                                     .readdata
		.fifo_q_1_out_waitrequest                                   (mm_interconnect_0_fifo_q_1_out_waitrequest),                   //                                                     .waitrequest
		.fifo_q_2_in_write                                          (mm_interconnect_0_fifo_q_2_in_write),                          //                                          fifo_q_2_in.write
		.fifo_q_2_in_writedata                                      (mm_interconnect_0_fifo_q_2_in_writedata),                      //                                                     .writedata
		.fifo_q_2_in_waitrequest                                    (mm_interconnect_0_fifo_q_2_in_waitrequest),                    //                                                     .waitrequest
		.fifo_q_2_in_csr_address                                    (mm_interconnect_0_fifo_q_2_in_csr_address),                    //                                      fifo_q_2_in_csr.address
		.fifo_q_2_in_csr_write                                      (mm_interconnect_0_fifo_q_2_in_csr_write),                      //                                                     .write
		.fifo_q_2_in_csr_read                                       (mm_interconnect_0_fifo_q_2_in_csr_read),                       //                                                     .read
		.fifo_q_2_in_csr_readdata                                   (mm_interconnect_0_fifo_q_2_in_csr_readdata),                   //                                                     .readdata
		.fifo_q_2_in_csr_writedata                                  (mm_interconnect_0_fifo_q_2_in_csr_writedata),                  //                                                     .writedata
		.fifo_q_2_out_read                                          (mm_interconnect_0_fifo_q_2_out_read),                          //                                         fifo_q_2_out.read
		.fifo_q_2_out_readdata                                      (mm_interconnect_0_fifo_q_2_out_readdata),                      //                                                     .readdata
		.fifo_q_2_out_waitrequest                                   (mm_interconnect_0_fifo_q_2_out_waitrequest),                   //                                                     .waitrequest
		.fifo_q_3_in_write                                          (mm_interconnect_0_fifo_q_3_in_write),                          //                                          fifo_q_3_in.write
		.fifo_q_3_in_writedata                                      (mm_interconnect_0_fifo_q_3_in_writedata),                      //                                                     .writedata
		.fifo_q_3_in_waitrequest                                    (mm_interconnect_0_fifo_q_3_in_waitrequest),                    //                                                     .waitrequest
		.fifo_q_3_in_csr_address                                    (mm_interconnect_0_fifo_q_3_in_csr_address),                    //                                      fifo_q_3_in_csr.address
		.fifo_q_3_in_csr_write                                      (mm_interconnect_0_fifo_q_3_in_csr_write),                      //                                                     .write
		.fifo_q_3_in_csr_read                                       (mm_interconnect_0_fifo_q_3_in_csr_read),                       //                                                     .read
		.fifo_q_3_in_csr_readdata                                   (mm_interconnect_0_fifo_q_3_in_csr_readdata),                   //                                                     .readdata
		.fifo_q_3_in_csr_writedata                                  (mm_interconnect_0_fifo_q_3_in_csr_writedata),                  //                                                     .writedata
		.fifo_q_3_out_read                                          (mm_interconnect_0_fifo_q_3_out_read),                          //                                         fifo_q_3_out.read
		.fifo_q_3_out_readdata                                      (mm_interconnect_0_fifo_q_3_out_readdata),                      //                                                     .readdata
		.fifo_q_3_out_waitrequest                                   (mm_interconnect_0_fifo_q_3_out_waitrequest),                   //                                                     .waitrequest
		.fifo_q_4_in_write                                          (mm_interconnect_0_fifo_q_4_in_write),                          //                                          fifo_q_4_in.write
		.fifo_q_4_in_writedata                                      (mm_interconnect_0_fifo_q_4_in_writedata),                      //                                                     .writedata
		.fifo_q_4_in_waitrequest                                    (mm_interconnect_0_fifo_q_4_in_waitrequest),                    //                                                     .waitrequest
		.fifo_q_4_in_csr_address                                    (mm_interconnect_0_fifo_q_4_in_csr_address),                    //                                      fifo_q_4_in_csr.address
		.fifo_q_4_in_csr_write                                      (mm_interconnect_0_fifo_q_4_in_csr_write),                      //                                                     .write
		.fifo_q_4_in_csr_read                                       (mm_interconnect_0_fifo_q_4_in_csr_read),                       //                                                     .read
		.fifo_q_4_in_csr_readdata                                   (mm_interconnect_0_fifo_q_4_in_csr_readdata),                   //                                                     .readdata
		.fifo_q_4_in_csr_writedata                                  (mm_interconnect_0_fifo_q_4_in_csr_writedata),                  //                                                     .writedata
		.fifo_q_4_out_read                                          (mm_interconnect_0_fifo_q_4_out_read),                          //                                         fifo_q_4_out.read
		.fifo_q_4_out_readdata                                      (mm_interconnect_0_fifo_q_4_out_readdata),                      //                                                     .readdata
		.fifo_q_4_out_waitrequest                                   (mm_interconnect_0_fifo_q_4_out_waitrequest),                   //                                                     .waitrequest
		.fifo_q_5_in_write                                          (mm_interconnect_0_fifo_q_5_in_write),                          //                                          fifo_q_5_in.write
		.fifo_q_5_in_writedata                                      (mm_interconnect_0_fifo_q_5_in_writedata),                      //                                                     .writedata
		.fifo_q_5_in_waitrequest                                    (mm_interconnect_0_fifo_q_5_in_waitrequest),                    //                                                     .waitrequest
		.fifo_q_5_in_csr_address                                    (mm_interconnect_0_fifo_q_5_in_csr_address),                    //                                      fifo_q_5_in_csr.address
		.fifo_q_5_in_csr_write                                      (mm_interconnect_0_fifo_q_5_in_csr_write),                      //                                                     .write
		.fifo_q_5_in_csr_read                                       (mm_interconnect_0_fifo_q_5_in_csr_read),                       //                                                     .read
		.fifo_q_5_in_csr_readdata                                   (mm_interconnect_0_fifo_q_5_in_csr_readdata),                   //                                                     .readdata
		.fifo_q_5_in_csr_writedata                                  (mm_interconnect_0_fifo_q_5_in_csr_writedata),                  //                                                     .writedata
		.fifo_q_5_out_read                                          (mm_interconnect_0_fifo_q_5_out_read),                          //                                         fifo_q_5_out.read
		.fifo_q_5_out_readdata                                      (mm_interconnect_0_fifo_q_5_out_readdata),                      //                                                     .readdata
		.fifo_q_5_out_waitrequest                                   (mm_interconnect_0_fifo_q_5_out_waitrequest),                   //                                                     .waitrequest
		.fifo_q_6_in_write                                          (mm_interconnect_0_fifo_q_6_in_write),                          //                                          fifo_q_6_in.write
		.fifo_q_6_in_writedata                                      (mm_interconnect_0_fifo_q_6_in_writedata),                      //                                                     .writedata
		.fifo_q_6_in_waitrequest                                    (mm_interconnect_0_fifo_q_6_in_waitrequest),                    //                                                     .waitrequest
		.fifo_q_6_in_csr_address                                    (mm_interconnect_0_fifo_q_6_in_csr_address),                    //                                      fifo_q_6_in_csr.address
		.fifo_q_6_in_csr_write                                      (mm_interconnect_0_fifo_q_6_in_csr_write),                      //                                                     .write
		.fifo_q_6_in_csr_read                                       (mm_interconnect_0_fifo_q_6_in_csr_read),                       //                                                     .read
		.fifo_q_6_in_csr_readdata                                   (mm_interconnect_0_fifo_q_6_in_csr_readdata),                   //                                                     .readdata
		.fifo_q_6_in_csr_writedata                                  (mm_interconnect_0_fifo_q_6_in_csr_writedata),                  //                                                     .writedata
		.fifo_q_6_out_read                                          (mm_interconnect_0_fifo_q_6_out_read),                          //                                         fifo_q_6_out.read
		.fifo_q_6_out_readdata                                      (mm_interconnect_0_fifo_q_6_out_readdata),                      //                                                     .readdata
		.fifo_q_6_out_waitrequest                                   (mm_interconnect_0_fifo_q_6_out_waitrequest),                   //                                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),        //                          jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),          //                                                     .write
		.jtag_uart_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),           //                                                     .read
		.jtag_uart_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),       //                                                     .readdata
		.jtag_uart_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),      //                                                     .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),    //                                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),     //                                                     .chipselect
		.jtag_uart_1f_avalon_jtag_slave_address                     (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_address),     //                       jtag_uart_1f_avalon_jtag_slave.address
		.jtag_uart_1f_avalon_jtag_slave_write                       (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_write),       //                                                     .write
		.jtag_uart_1f_avalon_jtag_slave_read                        (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_read),        //                                                     .read
		.jtag_uart_1f_avalon_jtag_slave_readdata                    (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_readdata),    //                                                     .readdata
		.jtag_uart_1f_avalon_jtag_slave_writedata                   (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_writedata),   //                                                     .writedata
		.jtag_uart_1f_avalon_jtag_slave_waitrequest                 (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_waitrequest), //                                                     .waitrequest
		.jtag_uart_1f_avalon_jtag_slave_chipselect                  (mm_interconnect_0_jtag_uart_1f_avalon_jtag_slave_chipselect),  //                                                     .chipselect
		.pll_pll_slave_address                                      (mm_interconnect_0_pll_pll_slave_address),                      //                                        pll_pll_slave.address
		.pll_pll_slave_write                                        (mm_interconnect_0_pll_pll_slave_write),                        //                                                     .write
		.pll_pll_slave_read                                         (mm_interconnect_0_pll_pll_slave_read),                         //                                                     .read
		.pll_pll_slave_readdata                                     (mm_interconnect_0_pll_pll_slave_readdata),                     //                                                     .readdata
		.pll_pll_slave_writedata                                    (mm_interconnect_0_pll_pll_slave_writedata),                    //                                                     .writedata
		.sdram_controller_s1_address                                (mm_interconnect_0_sdram_controller_s1_address),                //                                  sdram_controller_s1.address
		.sdram_controller_s1_write                                  (mm_interconnect_0_sdram_controller_s1_write),                  //                                                     .write
		.sdram_controller_s1_read                                   (mm_interconnect_0_sdram_controller_s1_read),                   //                                                     .read
		.sdram_controller_s1_readdata                               (mm_interconnect_0_sdram_controller_s1_readdata),               //                                                     .readdata
		.sdram_controller_s1_writedata                              (mm_interconnect_0_sdram_controller_s1_writedata),              //                                                     .writedata
		.sdram_controller_s1_byteenable                             (mm_interconnect_0_sdram_controller_s1_byteenable),             //                                                     .byteenable
		.sdram_controller_s1_readdatavalid                          (mm_interconnect_0_sdram_controller_s1_readdatavalid),          //                                                     .readdatavalid
		.sdram_controller_s1_waitrequest                            (mm_interconnect_0_sdram_controller_s1_waitrequest),            //                                                     .waitrequest
		.sdram_controller_s1_chipselect                             (mm_interconnect_0_sdram_controller_s1_chipselect),             //                                                     .chipselect
		.sys_id_control_slave_address                               (mm_interconnect_0_sys_id_control_slave_address),               //                                 sys_id_control_slave.address
		.sys_id_control_slave_readdata                              (mm_interconnect_0_sys_id_control_slave_readdata),              //                                                     .readdata
		.sysid_1f_control_slave_address                             (mm_interconnect_0_sysid_1f_control_slave_address),             //                               sysid_1f_control_slave.address
		.sysid_1f_control_slave_readdata                            (mm_interconnect_0_sysid_1f_control_slave_readdata),            //                                                     .readdata
		.timer_s1_address                                           (mm_interconnect_0_timer_s1_address),                           //                                             timer_s1.address
		.timer_s1_write                                             (mm_interconnect_0_timer_s1_write),                             //                                                     .write
		.timer_s1_readdata                                          (mm_interconnect_0_timer_s1_readdata),                          //                                                     .readdata
		.timer_s1_writedata                                         (mm_interconnect_0_timer_s1_writedata),                         //                                                     .writedata
		.timer_s1_chipselect                                        (mm_interconnect_0_timer_s1_chipselect),                        //                                                     .chipselect
		.timer_1f_s1_address                                        (mm_interconnect_0_timer_1f_s1_address),                        //                                          timer_1f_s1.address
		.timer_1f_s1_write                                          (mm_interconnect_0_timer_1f_s1_write),                          //                                                     .write
		.timer_1f_s1_readdata                                       (mm_interconnect_0_timer_1f_s1_readdata),                       //                                                     .readdata
		.timer_1f_s1_writedata                                      (mm_interconnect_0_timer_1f_s1_writedata),                      //                                                     .writedata
		.timer_1f_s1_chipselect                                     (mm_interconnect_0_timer_1f_s1_chipselect)                      //                                                     .chipselect
	);

	TOP_MSOC_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	TOP_MSOC_irq_mapper irq_mapper_001 (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_1f_irq_irq)                      //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_c0_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),          // reset_in1.reset
		.reset_in2      (cpu_1f_debug_reset_request_reset),       // reset_in2.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.reset_in2      (cpu_1f_debug_reset_request_reset),   // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
